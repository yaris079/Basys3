`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
dTJrc25R3smFJ3/BdSpCgVI7Do2i9P2SrWCjRFE2EndIQ9foQL6R358o5nu0gdwSq2jxocRZBvDo
WskDAMzOig==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
I/hWyl78NXFbc40vMsG+qer33YQM05zyiwz8/DtO/LvMqufZ/Ti4V0HTGVSX9kff4HvRLw66i8DF
HQWJ7R6T16JMIdVoX28d9sWc801kUMwnCvWddc8U5YsbJROm07xdOnCe6qWQx8GxZQjUTK2cIH9l
FUsr6RPrftfS6YMXxdY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jUGMkd4CCeSlaH93LC3J8ArSOZ2KVDjQqEu6hBIHvZsG1CpGqdquCYxRbz4ZyiRxSZ6iHRBz8BOu
h1ZWpCRnR1B/0/8KPs4Cs+cBY3ECvqp96A+Zd5NANddFRW5Vvdof9bigxMNJ5kz1phFjvUG+if7+
PIY5xkiW8/w0RQS97DpQcqgebLChp0aGET9QKoeSkrfwg+VHw1VB/9wtTaJd3+1H7YoE6Ullo5dn
sCH9A6D9pjjEkf1wswDVmOzq7rkV87nEWvx4+nQCPifBE5N7qMyD0VKv3vDE+t6YWoYFu08SRwf9
D9CZ3TY7mahKIEyiRbMNJDdafYlxulJOZhUt9Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jGaDwnxz/3UuoQw2sfeSH8LbEuopjExdzBLenAfAQ0IbFuwepeINPx+iFnbi0kP+EHyM1LLsMV9r
v/1WLaaYXLCcIxGk/7UKK5BJbgYPZtODBwsWBPtyXzalJFE1KPo6HEBklajD0wvFvFzo/4RLlzyi
cBhkjMYuPZZnfdzAC6g=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OMlubMGW0hm7AEM5gzOJHLw2vxYSaZxHswt2M1JGBpa7a/tjk+Z+8U2Qkl0s0HrPRNos8JvaO1Oj
xD6kCbPztsRxwg2e6gjqYC/ZMGZZ+oZ7lard+oZJe4XGlIKaXBjo3XGS7rm8KR10b0acOolPszRj
qjt8xp/T496ltVuSd5uVVT0ZC1UfUV4APjX+ZtlNDmvvZZdCaFGBDVBoqkMPZyTmyNJTPMskc6yI
oNROGEhhgid1yxaiZ1g03ZTnpc2+VyN7xASUXbNMm+vaYoPaZvwMNOw9ndph08ZTB08QWGkHe/ul
M3cAYfxOYYIo/gqcK/PqUBu40L58ORKWV6++tQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6640)
`protect data_block
K0pnidCqV1BarET6HPckOnQoNLjS5uW5JZkrA06tdpWwqk3tzlSQjkt9KAiR+gI9BYjzr9MS3QDf
BGJMP3BHRtSLTIgJ7UoJCRN5WiEmpBPiERdroVlIzyK8ZKfgoNjCCMX8H3vPhT8kMqI4YMB4OdJj
cMBRWIZTqZUcUJRjEpuuSMZqwnZ12aO41eiWSuuX8V7arENdRsxYGbkdHj3wwoJK7A1PHSjANInT
Z1X7WgWrWf+HuS8HGhrYiucLIoyf5l0G4A1kEqPROQTsNSdXEPew7tkWC3iHU7NeE0simuu4FQQc
xklV/csZ1TwVtW9lyuJaR7kmvlcc40UMub/IzW7f0X5WZqFOX3T1SgDLElZp3RG4skdJcLh523lw
juwPWDtAwwvoRN2cfX/PpZ1nlTd0qJOVmECVlDMC0Q7onJLgKAvFlih9Sr/OnsNeEeYPvnEEhQkK
dhZoRTiuuKGKxLEfR8n53XB56amLXE3BrHRBGy5CsTaoULCpTa/SSiNc+4lfh5Jr7Ij6lKR9SnGD
nXn/BMqy96uIFp9nNwbWv7uL9n2h+AC8SkKfygt6zPRPy4ZwEqprgReDi4kzLheHmBRyErVWDJuB
k8TqY6ydt0WtyLsuAt5VzRANBrINNCNBLxVjsHEcG49r6wrB4XfjwlKg/N1JVeE0bo2AIwtJB/7E
UrcaSseYfvgGCI3x6XQadswLEHpGEnRXJ2fI896iB8C+Zus+NIErvRgUXmqd2Nv4Jkv0ir6593YW
bySR0PLIrp+s6cAX9Pl06OgXWix6ZvzrIkjRLw4JcQIiJhkDfoVcTmi6pSfKYQ/svTONfKlU19PP
S2vbUDvlboYDuhl3Ca6xrojggApG+Do3vUJSGx0A1DXWLGj7bbuhEOSCIIICv/08q7cw1cp51hnG
AKK13hoAw3c+L/YAV5KOhurePv6w4pOMKJ13V2lzdD8e5hrJ5O8DfC5Uu+mGyBareAybgkVxysC+
EyVBll/YHRCP1qt01Ahd4cLTcUFLw6QFHsIntSZiw4jdDuW0sSVh5rkeYjuZGEGGJpJMsAQgJb3A
LB0jY4h4O5+g14sHBJlkPIHJk1N7jxQs/lyAeqHyTE5ZLemCfj0j03xTcGg70EiIg12njkYyWvO6
enghkkSOyRvsgw9L2np63yF/CT9K1EZRUnjLv5oo8jmLcsJedjiFXrBCyGi8LFrFNP/hw5tYfHTF
qzp19bfv6IyfFt0tJ2eQU6S+Z0Kyq1xu38U0Jxh+K4gMmbWgOMoVFCwBe/oDI3FkTjQcvwoy+yo6
cgf2sOd4ktQlm8S4x3HHv/UhgYUhsl7Vxxuhs4H/L9Ey+icq+dJcAEtwHASIibKXvVUv1RXjq7ly
ZSuPyGa253cr8v6C828+zSn1KEzgVitBupYIIkmVFB7dXJRt1jZmMjAOSrMisdBx66/iPIlmWusz
i7omKbwIkfFrzEGjvCFpufoD//Ax6rH1FENMw7Cr5FuRm4uXKhEKa7gWzfYdxdLeeKFrQt6g3zs9
Hf2f+I9xwIWHMe1z01WNkJGfLtEctQKQWD0aueaOMfWW1NfrFnny9oG38EpfNtQOAOg1sVBE2Ebk
jY/i1n7pAFSr/Gvzbwtsb/tVLDC+Uo1ov9hg2WEkV6ykMaxrgONNC1gELSkRcQKPJL1YccYhInI7
NGAtpVeginrPsYFYfZ19crIKk5IFOFGPN/D2WuEtZXj7k3oMCAuRmGO/vEZ5mlTzf1z/npzK4KhH
1dFWxXcniSfKUJI6ero4ozjo6gW5h+NDHNc57OKQyxpMgsZqu15DAp4Z7Y2RNDDSl4TAEXZ5+OkW
sSizG/6YUEcqu12tU1OVfV9lKk4oUU1xrvRVIL53fQgY1hkEevAG+TwMFa7ehMlPz80wP5WwORrU
m6nAHHO1pzsqjgQanV6+IvW29K1WAXJchEk4sFP4nbtFSgeN/wMSgBsGxJDCRvpQKCHooMtnpnsV
wpebv3DOSWmm6XiM6dNox/PZvXLeC28fPANM/fa4u7UqbiIOQgA9kfY327Lm89EiSf7alnMOPbVu
PuM9mLj4cUVT2pL8g9ZcMDyuuZIdHOU1BpgnCXNyFiuBBE02JmJWEDRnPlOG9qKEfz5NO7J5QHY5
S1O8jfXKZoytxiBxwxVXwZ+u7Xwuy52Mesz3XlVcAWh/tfgtSMM6EU4nrqId32sl13sLlkCljVzC
KMVYahtH9+qccSFfMrmTLoZ6hGMBpoJFmwX5HE/vVqU+BDIMeq1X+31B2IC2IPvul4O1uJfOcxhP
snOtt1dXK7ZevRGOXFgqLA8iA+wypunzzT/gX9ozoQeChiyFjK+RAuGROWXVAPuaxHyiMQFx2p1n
0boNvveEqi3I5Yx+lp0SIkXGC+j77LwxiyhEwDwXt8uQJcg8JqMhlSLBAaWk6eeyv8FvgKESeLtI
9BKy+LBu/11Y3Z8oG9D1ZmXmS1vDYBgSVPEGlPaq3Q2nZHg+E2L+Xr6qyF9f2cnlLF3zaC4M570e
tW15cF6wGKgefhB7CPLLFvHvTF8GmJYdbEHax7P/RB/o1XrqsAIUthPYbuzkg4bOHAxA+GZYisAR
bmnrEv5IVMOoqAim8DIUNORYEmros8QkiORvM0PwGleU0KBCm9Y68HNjeB1EQrxvQeDeZJakaYQx
Otb0N9uLOf0a28DCeaOu8yZEyR0BYsKIEGUCY7anbZzOiehUFTJgQ/jFOc+sbDboUsrMnAxr6v9w
iVLFbieEQ4885/Q6MiAJ/WGve9RHurLExPABBPTTbCBr4aag6r5vfXdV2bd2snB8kBeDXbrQOW8L
jjjgfFNj1TjQKRbd073TXtxWDBMaPC5O9rlgRJgSwmfiVbtyuqjIg4cpxSxKkM8567Fieogwhk0X
XQTxsWN84itzh4LvcRYbUUrzSQGI1o/6f1RXVGjkJOx6hyXwbQsP6CicUb4wW0ZVIrIkYtkD3v3i
kqvaV5JOpJhc3TgkHbgCv/SjtbFWRpQ3CXkbDeIILMea5Z7sD8sDE0VCY/BKGi+8Mx53aShaemLc
oOxjXiYJIfdGwVox84yWWJ7X/ksDC1mH1cnYR1rkzzH4LWTrfgexeWzNe0WO+lA28tikmSWAqZdY
YUiYatnFytWwpuyZuXtcGfjWJvy0lHYSQJyhb4hPF+SNiFcyeBihFTfOg8BBvCIrAA81Pd94F5/l
Q/LUv5uBVHsgdMWD5rOoPiIG4jK1v6Ri5NyGEfkW6ATnvvGa3jzJJlV9UuawkngsjwUdLMTy+tvC
qdG+NGQcHuaxGB+JN7+rlJzmaX8xSplPbCyW3ZJI9tEowfxU3zYl2xC+5FqH1VZmkuWSNJqQDjVT
/ekBm392RwrX0F7+zXI0FIUO1waffmPZA6kImWyLE+THPDhUn67we8JpiKjyjHZJ709kTwucmQx2
1IBVH2IH0o59G3wM/TaPso8aCOr7vASYhuOakdbusKj+os1swKjxicFfPcjnUmlI++M4Oh1wYR+Q
0Wtz/gM6yN6TDoyV8qej4GW0rwR17loTjaXUaVPAV66jKKgtVoBIq+cGR4/enMrx/UEVhz82tyZT
g1o6jzxtaArNml6jpae2hiSqTOHlFAqjtnDYHHt2XUTAuPfUs428KLZjcMkvxy7QD4YXOVvuVKEk
0XOjFGvmHnqurCfQCvgcZj/quCm5UbxS9MyK+8YC4NrtzkHnfN8rrO8rn0rv5mHat2F+yKmMefVh
t+CNez1Sj+12h/j7xwXE+4jGlB2Xe/gi+8q7Y6cYq/3Ki8hO3N6j9jjLxES39lS5Ez8B3v+qizsl
PWitGLjECes67WvSl1p4VeaQ+hGSNHiZ/Aq4si4ThuzOhjW1XwDe9UN14rzQwmj7dvhabVYOm9BT
Tu1gXmoGJJdvkChbx3AOdoQqEjIiRnm8+OvfQAI5QJGcsj5tEgiuG8x2U04igFJsjrBKXQ5vfLdI
DFkViL9mgtosNcTrQaEBTCjHDOAuxzWLEASBM8DLiLEawRdzshxSNuSFWrz6sZUAuVWeJUWMYtDA
8YRUieh50zWNbayfTpqh9+2LBb7KTmdyCXTUOi2CxQ4MIl63RtMWaSRLrblqsqn3/4yDmBJ1PDRU
XoQM3bRBVhFRvXb52u2hTovPvB+UbI/QMNewUWn+5zITtl/I47ZZzouFoThDnXhouYBq5cEg+oYs
5AJliHKZuzXqXq6VNBq8wb+kxuFyvouCivEHpPwMMFNoQUvMFTZ0Pneqprr8E2Qy4YbNKzBrEBjP
jLZ/HTVDK3ypKvCY82GDHfL9sKvtERrfKy/9cqCfCpAlKt2WSfJzFW5/56bduD3sai+vCCbPUrFY
ikrZFJJ6jH+yOkhKmugbp7piVNEM9AWni1bntwUIVe7Oj+jXoDZKGlNGtNFgUZEeu1Uc5MHWJ2f9
+hqCW8feQ0XRrS8EjyJ2tp0d/0wcHR+d9zjB1GLSB+k8sL1cP5cGNxvFbERbdsG9dkT7k9fbfpoY
t63cwEGe4J314+KxuIpST4CIWBv5TwBiOiNUbbfC/0eUffD88KZHQglvUm16IoTOo0LjftmvNOun
CG7lxLU10v60dUnCstuTqk1rbJ8FnAseudgjynnz3zFWXYm5IswPfTXsDtSqQNugvpf8J4ZjRO15
Ldket0+N9pF3zv9SVxv2q+UmwQzMTJ75uVpvytvmwY7m5Vald5oJxrlh+xRxG9/18vaTRcCjRL0l
JuDjZTpXXnaWCNEoVVCUswiRunjiFSRHFUdFbMEKRevsceV+ya/3Q3WwozYRK+VHSQgbC85lg7Kj
Bf/4ea0s8ZxPSpr7vZFlCHIR7dRGGeJ6yotOaLnQz1mCsi6NVzjVPQgypCeDldLaSsPqtouxfp3i
E3LiAWVO1b3LCZkKFEi8JJTVysPjHCBfyPC60Ow8hdJrW8soNdKYo12xFT0GAFFCb9KusB895uTL
PqoFoEj97S3DGoBBDQZ5rdzXRaj1tfxe9eaxXYoAxpcDQIElBOL76mXECcZ2Ll28nWbYk1fOditZ
+3QD+rtBsTj9RixMHSbyRLRuR1FJJPD5Sw0EmtbKDHCHLOwRRHzUDBzML9Ik+v4uLThft5zhAeJ5
OBznhy+4tKHt13RMw1L6rTFaq1ViBF30WnavzG31kzaZNUKQuyueFrP2MPzxwjSsCpmmwelwu/Cl
6k4rutzvyf/grb6mUQOubxde6bD8a57KovAft+BCVfhxL8g6QpiWpGrIfInD63sOmjwIym/k0uPo
M1FbNXjwh8B15xAMH2lHjbohlYrYIadggT+9OEx+j6xHvtckgitLumdhgB7InAmduX1BGzbBtGJ3
yjy9cX84Wi+2s5cLpeaRCIONhE7fo2Ctis5e7pDIqyISiYE8vzLxFN+glydyzfFgoid/trT4vDQL
QS46UIRulCN5kiIsgO+WuJh+xa10KzJCknDTgV/i/sCla/xzYKIty158Wrvdfa+rQ6rqChitgU/o
ne2hPkEoJE4DYV7FHAmr0zlnNvjGWmzsw1IHBUdZF/RXr0nLZ3Z///7jP3KH5W0+u8jQSkqy994j
cduwCnMIx4FUURh+mtumQLXkCRYH6Su0nCAm7pVsrriK1307DNz9dQqnUMpXdRyD1/PLdoW2sCzB
ecJWg28A3kspKzbTZu9W3PlczgiPZ7M4buF7/3qr1DaqESIxZD/xC637Me4vWBBJDtRSEzXfcIyK
M3xfbXjcsHqVSP6qj452VGOumngNbSryV53M7K82rgAfoP7+9+MKl7u77hLlIvqntPm/8Ns9yVGb
DwfI/2LlP/C6Rlk9/HY1UTAdsiBRtaroxalHjSiDRtXj5ycgt54jnLD0jVaN8hQmpB0eqGqKDYbK
VdRBaZWOm0i+zKxeSd+3e2X6Pp0d8AXWSEQdStQfntVkg0NcVKjGjPdQnhwfH0CIQk8AVwFZc0Fu
+9+eCPqVd8olj95ltQhnBsatOiVdhM8s5Lv58aCFDtyf9rcpGXm/GLGe2zZlYc8Q/lpjbrKBhI5g
bqCaQJFZzd72FVPtM06738ZXmJI/fnYuqYP3uinpe6LgkYVgG02KjlEAoqVsqU5BOrTORzxp4ui7
Mx95awtGCQXjM4LbciTZR/EaN2rUGYOTDn58RQotkyqmUyvmsMvxbv1j21KpXgmoqEXb2M62JKYz
dvXeqDLBcAfeSvr3Y6ZiB55XHy3MWNDrkw9l6JvIBgPGFmx6vKtVytJbDqoKSIQmraLY1LuPC1Ml
ZRaQb4vpdSAb86Ija9tnW5gIHMPD4kSr1qe4Kd7vTHe8U8QzyTcL/UA7zp1+5cO3Wiji7G0IzRdT
m9+M+3dMM3aVm7U9IQVoJUUBCeuvus2cG1E3lxs+8r3p3nNRhNXJ/LhTVdLTimEJA0+23FtchhuM
qlJ4lpHOpRG5Sn5dQkJdjGKv6O9y7PFVEk+arW4cFs6rQPbxHw1FUk6n5zUO1oxXdrcZQHq6+mTr
9omEGLPgXkLJssaybp7aythGOSR3SMI2GWAMxDNMGGe8+fVX5QzP4l1y4v4UCGFgUTf28GUIQwuL
m00AiyUejvDQHin11gZICUU+bDwW82odM4EgEGf9JA3g4RTTX3CdJpMIT/UnT1jY49+lcXmV/Max
XJR/Fid/Se7cuR1Elwa2W0zy/ysUwiJu8yuFnZ0mzlV8N3VUh8PkeVcSnvzEjxZcPG9fDsL4peCK
Vjdk75NaAKGraz7TXdh+cpmbrka8FCHY1BCnVThOpqqXwYA5CyFDEkBVsVg+5/UcjDNeBJQGk6jm
8VBsUEKbnjLH2zmzsRFfpkwYOYQ4nDogyjeh+tMpEuk53KBvs1rzIRI2V4sucjPKouWpX7qiuLRN
KHYxxWbsVwjh/f1SXM21XHuIjL2QMV67qU3/QrFPs0Kfv8+mLaz7a0avXlKJoKDD9tz3J/u2PytD
/z+RT+jsC5ZxLU4tz++i87lEL929g4uIT6og3j3B/awgmN83LFLGTvYnFnMWVIrqUnp+Sf3ad8/6
Mj4WkI8klUphTH4PnTCvwgrjD81WvWgfxwQccl5BfJH4OQ35VHVPs8yI2Mttm6cgZduTZjS+OPDa
ggnUP0HOCxBm7r4t1ggwqrHrMb2mnsDbqZ3eK5Xu1Ymt4SWr2IwvhgbiJis2b51oim8RjrQFVAnz
gCZGW+NWixcdFa05uaZxXpSeV6LlEmAMxoZKvExz25NMVfRYxSvcISsiess19RJ3Guca1eNfL9mt
HLpphXIYB5dC9YbeAGHzPY2Lepg4IjBjSnO8XbjJmWrR1WZaHUkLxxiGLB5w5PrhTHSk+RX0Xlus
XkqfjRd7TuNVdGbTUvb6WE+NOhM4oA6B7xFDKLvn274fEGfdn+VAPJB2k/EcHmniHpTjDEg53Boy
cfkytQs0tnmW4IYFVbxP1ywe4qLYSVf7Qlt3J7mGSNdNYyoqT4vmyU1H1RlvLRyHcSQyMK2TKaZB
Kug3C168RV447faCsPLplDAMLja10dm/nYG8/vO1TBOpEIwv55TCiO2uwzGIqGJg60tS6oG8DxVX
Akj2AF7fh3QZsFvbIxnA3jLhVG5etETYOvUo2fwVnPD3jJFtrqGIUzPiApctbiSx1ll6trpt9eeI
CVLOARaHWDdsPWLCmEBAaZbfJx799n+2BzzjbCgqrfK0l0O3Ca/oA5TUwe9fKxsv8jDdJwGsvCgz
2Y+9pCljMbO2RKIAdNUn9WWUpNj47RiB490RJ25W6Wtvz1w7konJnAsYfRownVyZoeqg+iJidNQi
Ai3JnWCEVuUzmOIct4ZvwPfKuGT00I/ZzryOeTwate0xeXnXjDHIPO1Cc6Ysr3ANjzuPDIVlLNsJ
NcKEr2W4DvdXW2XFZ2Nfpi4WgkCv2l4eCkKHmIKRa8lm/HnKiwUSLpKPlQFkd88JdYmZyVZGF1Kv
5bfzLsK8sNsmNFhXD8xRv73HxurxKc9m84EFfS+WjVWrkYv/KPu7RMAPnRpxanwoTOGqJ4jN7ugT
gCk1A5d0pc5wwlAmBk1o6TjC0POb6O0Yt6I5ek2/pqWy1y2pVTmxkBJkqSZWIuNrzURnz89lluOq
AhWgHWgZGaVVqANhY/iGrV6R4copzqwcM1vsHFYmmD2S1XbeZabnR1Yf7tm0mr8IxcoDomMUjPJ8
llmgUIJlOefR6EGBEqwWy3vBGJsg5E4LSq1y3KtK9lwDZsLQ7wBoaBI3SwFzl/3InqSsHK3dDVfE
9EyC7yijfrJDF5pe+chjChcimVGH+OHo/PR1qe55zT7PoGAJGaoFUIie+TtXCRQWUl0moxZ0wONy
Q1fFns4mYIgCGBvtWMIXQDMIDkTOEKb2XE+Kpb/v4UGXKJ003GlhnkuGr4dAMpj4f4+4Ld6uL9yN
+44SZwR+Ncl9PrCRvV77dpwTpZvzzpKP8+53obdiawXxLYQ/AYMJyeU98ZfMU8TcbDcrHzkRIYBX
XwaYVTy4oK24bcRwR8uvTbkYAcRdhjp091HIYnLpAmuqJUvfYcR5ZrrmlyGbDHPTcuueOqENn1wq
S7gr77DnNKQ5apwqS+T2XN2bVdHZbvayfI9avsT8r3KroZDuVQ9LyRwlBEeWjxEaZa81KQd6IhIF
j3fPy/rtIIGvlfERgKv5eFAr7cR2meVn1tEUtPxm9gh5+KaKiKYAnR9zHIkbRuyyn1DmAqqIp6tn
FZDCvg6RXXNf0Gm7zyT6chXkj5Za8EudrffDSh46aZ78VM+f/dBoOCNLidI6zTstAwHtN5Kn1mj0
AdVHw3im+s3UNGN4ss3TMv/wCIsLCyLww8T6Vt6yRsp90ykf+ML0qfc59pYlO3b/yzU9yUSmRTBj
IjqJm9tZA1XOxEVcwZmoSNwOMJD/eRC5DMMj7g==
`protect end_protected
