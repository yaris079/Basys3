`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
kqKY015M0AguD340wtFmn2T4Wqd6uyV1XCbeIylDG2Dyr4e/zUXXK/NVkW6QtUOP/s7dX4hc/YVB
P2YxgP6khw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LHrIthoEUHUZ8ONIKRkF6J+d8PQiIn6+n978Kq466I134pqnc4EMiRkTkNFZtDc0JLpc4x+aOq5p
TnkY3IBPKn1cdLCkOs1Upqa+k2mAgvfYvPgIZTrXuRvnzieQTtKc1aYuaLQCNg71DtbC8aYGP+tP
KOKtde7VGeFNWceRb4s=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mehVKOXMulCt/akQMKvmpAmwd6zOXI0sHjBFiz1/6kKBIyTNotX5WN6BrGks8YxUPjQHEmaYB7LO
ZXsWujUuzQTLAgZJxMMisYyxU4mg7wHYMwIi+2IKRHoZdaqHlT3lD2UIyYEYkbP2P8ZaIQHceZ0E
mLBgeCy3KKtxSlRpOQJCilIoAZyYuqF9GCxBjFROu9x7bt7bCDe37Xm1acwA/oERUYgnaR1kkt5j
Gk57JD8PAs+Y7pQaGFFWOm3KnC0fm5K5AxYO5N3av4qPxP4r0nYJD9glSXDBJjpJ8q+44J0Hnh/n
71Ro/x7SkZJExxFuYJFOH3UrV8+chsJTL995HQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CtBUFH74EmMGY/yYcic8SXodoCCpa3E7afYNwnD3Z33gy/S+FPjmY2lMrZ0e38F4fj4IltprDYOQ
wfXk8I2HV9ejVzbTEfJp3AxNeEtZ1rNKTol+Esyc3W3fFJbqTq+uL3z++L73fzKqkMCTA7HKgebC
ZSGn5TbLkNlRgP4H1sk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M5qgnRb00n2zxk/SSGoLcvwpOOvvO0IaUHbiQb3U6oljahzxrpAqWAgujdEtpcO8DaqxOI4SSbQ3
GjIfGd03ItG3aHvugYKEHZ37GkZ+Sn9+D3rkWmETLUeQX637kXhyrrPelmitPTs2faaIlE1wuaeE
W6UFbcKPI9rfcv3qCU4zSZMUp9k2iNaW6+m55bs7XMgHY+7SU9AdPa+YkLck0I1ougVTRfdjmjQk
UMfmGuYtl3ne77MGjREgLIg13Q+AkH67GR0g4Qu3Y930JPRd8RH1GKI+pPF4jMvQy9bBzRleAhdx
k5iu6/7nH1jwjVjvxaslAu4vb+mx32rPrrW2dA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4960)
`protect data_block
L368nUy3LpyZzIkuSo4KR1c+Ej8k0yT2oSquvh6bcjCFOSq60XAK0e75nT6ujiBkiVqr/FvcLM3h
JI5uL0mb73AhHy946wj/JsO3jV0KNK1dTIlNkk3bkvFQ2uJQO+LyxEPnafmPR6bxim1caRdQkfo2
3CK7UulHMMDBvUCxySDwGWC1FfETXBy5nyHwrxZjE26hqXZ7beGv5fiEL+VOV2JodTmuvRWGy/uY
S5wb+mG82RGVXM8ZTiayRqQFaHu2hYqQ5ppISVw059g9l/XfteLQvNPzwVTDbZmO1d6C9OdTf6vI
LBFIl8bECOyAIZfbcHV/q78I2fIBBRgDvpvflfqneeLfOyrj44EQW9vzwVYqhwCgSuYHZNA08LNd
kOOApD7W/wXqX3qls5nERHtmycc6pwmYKmTs8YNR3e6W9yIqTJTxz4exsoF2RpBOafZShbRPEwIR
SQUmO65XyZyadTr3iK12Y4nGyu2sbaNJNVZCnzqJklposbXKbZiy6S5/rFz9ACHFL6kxXtiuPlzC
zKGAuMGaO4OPy8fBWH2F3R0aO7DALBy/bDfUtz1OSZ9uyYvz2EkgsgzxMkZPqNjRysJf6jOwu98d
wtiBaTvk0S1UB5sVTnPTzJ8rl9lpX8CjcJ8s1v970SFtKmhGlainT32/laD+jv4XPmHXD1qV3LXq
qg4j5crbS9IDZUW+FQzdGzSa8vDTagZZB+nScqEiVYo/rzBSFrEbuu++VCD3kQwMb31jFr4suqkP
jG9UCDvYr8E7U/wpTyCO7uz02UQsdbISY+GC0Bp4VgJhd/y+m8xCHxvvkWs9SJOguj3YsFEDLRYZ
zHOFOKaYCFbfFIVKzw3S12m3htOeJLjPVJoXsT7cibf88wFh0SE5qmjmUAZluyhXMYtpdqZkww9c
ClX0a4MjXQqv09RrBRd6CdVbQ85c7nfjOpWslP7cVpfM7Cqt4UTLnEJKPssOQAjfIWBX4Cmh3Vq3
aUEDg3LguD98qznr0a9jP6UCXUCKBHUuKGJoLolhsoihfceG/TWC46B6zpdMGSjz3IC9812nL3Cx
E+WPOzYVEvmKYMVfnpjWFYjhJl9I3w1geYWyWGfMNpEDVWz3TxyCS4xCm1IJwEw+038nDqirKB1U
LQCVLvhp1J+1LnR6grqjmQxBPi94cmUkFbwzVFjKz/C6kcCVjrBLgYC0MXnylGx+eakBL0Umhc22
6g0wsq7whRaB89Lr1bmr1KYfAz9cuH/lowehJLP8y4yuWieQkd8nv5T4NzFXOH+LwNixbMkM8gM8
jvVP4xBfYRMvkwHAU+1ihY0mlsFsFltyw8EQSZpg+VA9/eRn53VU7ynWkqpAmcM0pnbs2bQ+tYlK
JFf/rPrANg+/6lpDsD92eEN/P8E+3Pzj0GuG4bQIqGiR8E/Aj2i5TOp4kPDhWz1GE35HTeQhEbgg
qgpOgxLUE5c9snW7q1F3g6ZwZT9cBWN3qoqFs9fTx+UE4XQrmcwKimtgka7HYZS8AxxFlG43PR0n
bMqHb+Sib9BWwM+a58uN1gnbeIKDSVhbZEi5DfXSNb3dGuKAIB+bnrSwbJsS8lbeqkWoVd4Zrl6V
YF9uU+tGZiBgezAl8mUPEHAvkn8zrz/OXmBbov8oJiig9sKjj7SvxhouqYUJa4hpo1n+bs0ZCRgC
7YWqriUe6kEC1N3SzIW2m7ZVnExQs2mSitCN1cjMRxhvXdAzZlI+y5UzTFUEsbSDDXTFb54OOVY5
R5O53Gsm0Ax7CydMcuXAHYMhfYCkkH05CAnwU5uSMonQNflQ07plMw+hcJTZVxILvAR+Aztma1IP
kBmJ6GYtO+4E+vs4MlZfwRMUoV3CpMWS56y6zv5R6kARXBtV/kXVnUD0sPXMCcvXy6vByew/hYrn
v8t2sSA5LOL2OwSmyfp3E6qTo14Unb6g77ir+/oSLrP6FOFyJIC0Go27b3JYbHy63nkGcZoEPgZw
i5S1V+qwk8a+G624+g5KxLKlPOnS9jfC/mOatqj/sbqoq492AqIc80sXpL7bjtsR42PnIuhuM6+D
kxeveorkkaPm7wjXFKAgFb0ukqju9gUjaPK5CSMM6Fqw1k16/6IM2YuAOtXE+v3KHA2u5K/gx0UM
IFrzIuqVyZb9IpaP4DDf3NYikYg6OgmANY5Z2SXlog3ru9cN5tAo7tFZQWWxvaTHcpYmYGSM/wje
fxLzKGfI03lKToGMt8hUDPZbU1kWxR4flW5rD/VsXBseQKrtVeHc1oITKNxcZo/Pw/CzC+shWM+Q
fV2+YP8rRZkE5Zg+mjkTOqHTfQ5eZbNBH39QLZf32Du8+vlRJSuiUAR7tfFi2vNosODahcMWG42j
LpIeh+dlx3NGDgMt3/OMRtsY512L8LM9g2QgyfWY69cD6j05My553ZWw0TZChr12L0IQi2FIRz7K
XqbwA/J3sK0K08WzqdKAgEUbkKjdUY1a0PZoikhpLs7DvO/u+gscLivsVO6jXBA51irubDWhsWCL
xo9IFlov6uTgJrLHNcFDAPX5dLFyQb90tBE4k/jVn+2LwKOkZcyWeEZRf03tqzPVL37E1ofRbo1v
GY/B9hjunv3YTZTZ1rMR1fRuexvo88uhAr1D4/tsSizk2IoF1Gw7jMjvnUjduPQLPlYdPA7DV9cH
flIcIyCh6pToXb3ukVEE1FIbXn/+zp2210dmj3s/m1YFEgqIkap5TelNL8FLoKvulEarHG0iAhP2
xjjoiFEZvrabYJOyTwHf5M6gonpC49KYAaHTOHGb282yhPFBZjKGDOxldMlV0cqGS9MPeMghqf0w
HTwQ2hGRMGzqoW0FpNqNTtcmmGO0hF3jp6Ep7FJ+fYtA9h/wY6E2fNbYsY4Gj5WEO8Zfy/aqyO2b
OEnPllP1a+QveZQQq7J7/kGANYubYBXqjk9OxXtWPXZki8WKb64M7QEB6etTEdBioC772pKCV5tj
ZSihiXWq1u4hRNJ5z60Gu3QvXh+PEYP/FwN+yLM9I5chQ15MYKsP0iSrFuL+BfaFFLbTD9fb1KQI
8h8GPt43Izl9uFRK5k4T/GSg+ce1BrJ60Vall+qDzz+A9hDDy7L8eMrQRkMcr8QY2MjoGRxXObWc
A8uVqF8O2ZBuwt07ZWMwgHMCggzoaZuHQ6U8j357fuBiPnCpvN6LIzGBLA2GsmkmYaj1Orin5f2s
WWvuMAylBy7ghGPr33YVSoIvui/e0/+wC3mq+8z/Y2LahnF0SOTcwAMl+GXmLztlzoqY0hSaL6Kq
mD6mMzqpQENVrZymZPYwGOU8DSk4/EFjMtEMH0eD6cQNTk1KWVtDC+kiyDZJ5tz1Qh/hgaAlbvQB
QeGN7DLfu+rUA4Igw+GQOlMktY0QpSA24ZFoRmeK7bHxdT+FMNzPjJkKBHX9arllmpSYw/b2nxgx
r5/70FHVcPuIvcQvh3v8dz9oY0ZcpjSMZBhZkQYJB09/0nYGliPxcxQdfvpfOdihFunuZ+Nn7ZoV
n5w/0PiLpxanoxyNTBNmBzqd5CLXXschMJ4tAzkYweUYY66rvdldvqurnpB6bHF+2p1rsn+W6yA8
PKz6G2K9bDs/MZpg84f3gFNbdHBZte4dvzmc71CpbN1j0j4sQQ7UwaOuEbyJ7gDui47uaISyYuct
yQXwzfAbuOjbFz00jcxEcICuhJ7T8RSajV+fzjbnzCx6NLmiE+EGLm+mVx20w4IRRBxyCe2HZNgJ
JJY6KzXbSa0Y0kP4QpKDdvV0vpI/johnu8MfEyS1soS8MkMwlK8Y9Oj4Gw0VjGmfkEakOrG+xwvG
j93TkBC9Tc0ukGZJ99DstwHbkxw3esI6m26AUMLF7VAlVh1aqcBpedu3o8S4plRQ+vKZDTS1+et8
p4998Orfm630sglsEiTjTYPWbphCHLA6bmmfFXg+SjfAUmDF7xqdYv5nY73APexGX51jvQujOSpP
xcrRwZG216VcHTjLi4wL71AqonDafnhrzs0vtx6TenaCtGTlX84v7C22RGiaSr0piFltl4BN8Svm
xInx0PNJWOzY+jGLYOpaRUIFjdLhFhSIEMlNoVpL3tY2V9G19wVFhKVGCCC2g5bejkxulq3V12Fl
TmWMt6aBXA8GIlanCpLuXEoKh0vYMXYPT/dIKU9g1i9W1W4VdIPT7g6TrVntJix8a7zbLEKtkoxy
GIhZR8lBDnnfkNoXJycaYTAhW0Zz5fGtOT9qGEbUaFyMxCWkIm3JFlprtYPbubgSuxfZCkhmksq/
vwJU4R4YwUZaub8Lwhj3S/08xe7c7bLIBq9ErfqM63jaHPuvX86ifEnsT8yK13hVb82nTAXIGSuz
1Iy/hJUyYWmbZud557H7Bi7RCuSEcn/FGh1yEngVNfg0j0icOOVvBCL6hs0Z09eJs0CHU+2lnTm1
ONqk+i8pzB2PJGKhSqp7q7RYG2eTGvvjkhR/erSkRm953WhiEAqb2AAI9npTWL6/G4LCqgmy4ERE
3JVKDIVnhUmF6I101JlPO1mVXEllpfhLFCmDy3lgxn3Y4FS1LJxslwscz2azP22jkYoVeHqURQ7b
JbL3Yhcdhe7ribEBSY3QrWvs6Ktawbg1h/u5W4g7a1PFs32xFUJAOVcA+VOBVx5WTBpjWx/tdWn/
WpMK51g6ZuHlA2u08FITIxMkBHL8osZLgIK6NWquntCo3hDFGmT7ZjG7/CVJ6qP2tVUcytGdxKas
JNFclDY90iWKaWEw0TrdjnO/RARwl8GDfSfdTEaV237fZQsX4YI7md9jlf9jIlCs7gFPh2emW2db
r93FSLNOWckZV4Sz3hdivDTAbJMad4+OPobX9Pk+3Ng75DDrxfhNdsDmyk4lOM+BQqDs/6LpvPn0
NnPW6Yc3eT4C2Z9J7gka4rf5GRokcQmMy8Pkqg1ZZ29xrEPVXJ6fMPHm4LQuMfOIoss5dJE+FMUP
JjyonOLNTVJuspq1Gi096RlxxuCb7+tUMEcLE9PZa3jhNQdcQUfNbB9D18FCnOu8FiF8hOjaxiN4
vz9GEv8xeKtygeDmjYuCJrRe2D5/2PASyRrGKb+hL5m/DHSyLEYnXV7F9LORoCmJJ5L572iEH2Rk
jZZn6YAXdWKnTAXmQMKLxa9Kg9ULx53Q1Y6FQRPoYA9oFGvWZC3E+Dl1eI5y0x6wB3OAySFcdaJH
vPRIj7LDKKLhStnKVOoBeApVa6OCxE/ia87H4oML5JGEwOPtKmA+ZlqB147seYWWW5DjU0bYkRYn
OdgAyhYD+hMwjRnCqG7Ik5tkuqcI88+H+qFuNhVoj8YrwEgvTW18LgeNBMcjX3dXcMy3cF9xPzD9
fgsRcfHSTqJv2vV/XlptMihkVx8oB/HVZyQY7XXOiHVavrPePRAQ6kyQhIX/z2ydMqaoItzfr87H
E9XNd2khq2bLNZQcKvEzaK+lSRmgwcD792MjPir5ugMJpDec6BRTJVEWFQwadlv//3mFwyIAMost
A4BvRNkeFOKUgPw/xhRh4AQ9iZlsl3FxXf+vLUFH/Rx6Wsof1mZ4plz3t8M6he1A2taR2yZ6WPnm
TBU8hrgX6aMB2j5EF5o2oDhWfL6MAgykebimnXiTwqeBM+BS4mVvwW6sTZuBr7S6G3rsVgfGR0Ao
8/gEUvIKYi8woRt9iMktYHcnM3Qd9VTA0EB4xgSZmLJlh5KlpteimH11bQT2ADKQRjTNRVsZ8XTW
OZuih3+L3TvpA0Jcuv0NRDV8tf8v+jXm0sXJGFV6TI4N7pVGmwnHDJ98U+pYD8aX/Pf/24nV6DkG
z50WA2IE0RzmskJFCoiKmg/jN3CfaS+9/dSj6+Y1Q88ibUxVC1a+My851pcjDLdPlQ2HHgy+nTVw
4bDIK7ptYtSydi/s+lYVHJvUU46xnW/hyuSSA6NPfX+yF7tiXq4tB2QpFJhYQbkmtN86hDLte8Pt
bxoHv9rAt8fTfwunEnQySWSYsfIdew6g1AWErB0s+ywiDfM7yXy7q8owPLWMpteV3L1QYq64Np8x
4XEuuSWjhAmeQ57z0FPqLTlHWjsRQWDto3H2ESfcoVyJyAcLLWWPEyiNM1skdZBTWMulyNDWbigz
D/SeD7mE09rx0sMP8gmNuKb7Hiw4V+kBA2cFGCGR6nuHGqDaLx9MQVEmOE2eLyXHnjDWuU3A/39v
QzGlOZDWw7x4V+fiA/HJFGEGfI2YM3XVyPzktx9IMT6GRRriWYFoqlWXknrNERSuWWG12E/9Bg5M
/V/gHk13O0itxlRf2eEYojOgjIcKIavE7QoojWlMos7YJre494MNXd/tNv6OQc4doHNvuYnUCBcY
GF6nEiXOFrue7XB5lj0FGgzffi4XM+Mmemj6U644YDeuLgC8PCfNuuybr/0yWwkFxFqF8sR0hJpZ
MCtzCorI+PTNErgLgvFnD1jSZu/B2yaZK/DQ0xKZF+souxyAUjYHqQ3srUikBCDxoQrNB/XbCzUg
cO4S+dJTGKHWSQgbMwGLgVuya2iM4/eEK7Vrp32h1qOXJsIa/E+9p3qRa7vnQ7LjcjireUn1zkWG
v3QZPX/TN4rpKz830PH0k5xPPCcD7B3MjJNzXTVXlE3MSx84gwTPnMescLwAldHfULzhELQXZdXa
Lw==
`protect end_protected
