`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
P/PJQr1VNSWxEG5drlp2PQZ4L1Kay8RlIgNUgGJoHBawjc70hgM0nKGVU7NsOlNOzYLjm3xUdE7+
zO5J1RUAzw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Yi1FQ6CniIUGmUmOx9C7KRueonFH1bbz6cagJDPdzTE/EPjrwckJ1CXVDqWTnnMM/syZPHAXk8Yc
f6WnXzHAA4TrCyxha3mhwN78Nfg6IB4rcNVsONRE8re5bncwu3Uo869fDG7la7T8P2jTxDsuylMS
pURTsBf2LG0czWb1SBI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZVBP+29EpNGwXdPswRW0s+AcW9BREbFjdU+8AY6pd4MQ89jrvo8yIhSuG+SZCTcj0epSBsBYSmct
75mor6wh1sYujIOH8uDRnzgDguTQFfrq/iBQGQ+q7jiV66+CpuUloQU5YbyYkP8oDhbyQAqKIIH/
eX0rSpVHCvKvSU615sfM4Rd6A+cX+2SItlVhuYIiMjHtfLjxZOOil5+XoKTueluQXdgnRgd0QyQp
CyW0CbhHFtH0SCn/c6VR5TgVdvX0b71Opjq84bl0C0+x2E3JbK72+Jd8A7JMgLGLYr2tMoa5Imdg
memX8uiBqlEjCAo93eQn1LVXUPZPMe7plzNJUQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QswrPUW9nhGrLibJzVD6XFeHtnv8HzfB+4A9rR7Pw7hcu1OSbyAkCGZMXaMXhwFgrQE/zSInO24j
UTYk98o74oavqRgq2ad1D8kD2RmW/vmldtlOwmZ5yYCoyeqCBgohT6/2q0JKltjkjcpzILf+j9mT
er1E3jHX7Ou3kHUzVJg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pPwioWXBw0fsGDWGmlHzIGa5dUOcLVVm4Tl4tihcr66jpMHY20w76hqgBAaMUgNAv/OqWetQWHDr
z6fwCpSrDOmnuLLOy+ctmjn8/d+apK+qaiefOoqDfzBf639QEise05NEauz/HCVMqNggJVubbiN3
AorKYN5l5WqXjOXwEl0WsNZllVKPMxuhlgYMJwkJl39A3GcImEcmb6ah0YFYUKfoS2IkyROY9axS
cn6JLiAqmwo1gJXmnMkU2l+9J0y+qEn8zGYUuv8W/rtJmt8BfPhe9s3U13aM9Av4uVUUQbXJB/Ov
hmDf1/hUl2ErG0hai5XxYiWBhXLYPANvCEhcIw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38304)
`protect data_block
Rjnr2GRWJHxrd7bkqOiIgCsV2QGFOHiOhY+A2TqLfoHipKpgh0swWdOZ52qDV2CTzw7LVKLEL5vB
iV09jGyvAYRySqunfT9PjliAjcJSVksR4VxzCyjpOskGcgKHS96Ddl/d5cQHSG5FoSdWqQTO8cNT
RFRPVBuFBfQU+BGAg2lfxN4TmeaL5UP9uwnEdYUvrZk17EbhliVttMD0avKzDDxoTjAApJJqT20u
TbOqftoHvMNbX/FQj9xV6JcJJUljyDScWOeLrLTOxQQxVY7MPzU7G2tvC5hw9PZSWoL4jDo9xWRc
+rPLKgjVlCP3q1HZMZfzXRn65ou3ijzSBGJmQYC7LGyVC+nBWm+IuCY85EQV6xhUH1owmYW5ZMa/
+E9zJY8ocjzbq1XsPTeoSGRQXDfScAjTnpWfiZbnPmBlmOXYwYB2t/NgZPj9Qf8pUyFXs1ElBBqh
SBjbslBXNIz3kfpnIUcGKbLXqgmr/eyT0tqssfEB24x1VM49XYZo8UqaLRYJ+EilFieRqoudeiO6
ApfCkJW4CK7hq4wm0uLHUaJqq+t52QZrXJm9XKAEX1eEsuzGW8t8Ry+cn16oPWHtGIt39QdZfmwc
CCwv3AVlfKKcKoYB/D+c+fv0d+Rr8fPDAwDpStD/ezrYhsXchBcWX2pJo3GG9m1WaQUp+lvl4Wt/
KyXU23wKaaqJ4DCGCIkX0IW/cMh5c1cE7L+ROAdyP+nAdBlHWFvrLdCMaS+Tr1tWmeImnYNWjHB4
VtiE1atA9CKk+WDz3aStaY0X4A8Fr0Cp2hM2HplqFybwBFRbPDGhoOdu2OSUMoxsgSxEV5y9QQc1
w6sVTaTeLIY/V8nyTQgVi2lx2WGEpBN+/PqivZanCG13zQ9cxuFk9kew2/tEXTu8mspUO2B1DkZ/
CSPevjNGUCQbFkgNt/DVlIRGhcsk9nbp+CnjI2T1MWLyrRL+cm0gmAkVNqj2yHMtKyVbfFRu+g+I
91DuNwZ0oD3y85IcvverB+6woRpz6+aHuzd7LZKDzN5dSdxwjB5+p//jnfhGfSZmYF1IzHtkfxpS
31QGDX+jiVZsrUile9lxYshZsrjr//s9/Nz7dBHq9n1JeIzLpJ1bBZdJWJF+T2ju4jC+xENsP6Ce
zUQnszuSKKftkyfADjZjh/DpJAMlODN7zLfFO5TQN6VU04mJ7QW+0OTRZCukiaKTJCUv9+QszEJl
Y46Gm+JIs7/iZFaiz/OUW3oh+XjJa5IaC4lvyPmteOKhfMi1azmenUva7Ia7JbCKviIEwUksFYql
rcurXqUmqIIovYxL8KUH+5B1vHix/KL/AGk15ZFBCugQUFqHrhNNMNcA24jK1I2AtBX0wCWO+plL
fiHKDxoqdHKYzghzLBujiyLY/aq1F+J02FevO1tcaCot5pLRfVfXpJnyv4mQYJ7QaU6W8n9LUeQj
S9ADHPd9N8Vm9pQjYcNuwaj4rpCJmfel3aThwlgPkj9bEufkCCl5nTa3/oZsRj/4a3EiBKw1Zv9j
YAK4RGhAdxGH+jCtRa94AKCKOCjk/NMpn0D4Lsq2b74xKh2bzuMMPqzMQWT1OmOA6aanBeVkU0da
dDrCburqtHZi/NMkcnLORDRoZPRDLKT4YxoyLU0qKtCIbKlrynnzTgNitaSXboQhhkTsMpLi2FsM
1fC3Rr7HB5JztHuc54VUdz/lLW19c8WOVtz25NgRzSW8+6Jhpfde3FQGvpLmcbbtfZzXAblVWtLN
fPBqV9Nsx1V0oRoLNnX+tPfJX7vejSOC2Wk2Ai+J+z3qVK8QlAVEjBf4qbpqjnM5Kv00SbU+UW4Z
Gqea1Wcux6iKkMIiwB1I03+QPPpjjD4RwpBTa5PcnYjGRNokc7z+9+sMSAmcATrnUMO2i8OI+c86
Ah7PgDHYrUVFxpD3d7jkzG+VJuiM81yhkyCN4saWtA3das8N8CopaeBLBDR0YPXUtHU4bizPNmoZ
EkKP+970X9foz1doiDtO1K4djitOn7oum1q4CUqVQeMT7rpqeziClRxhOVfRU8AppNEpU3M8wfsl
RIqiY2cGqZIc8+f9z0E/uVfNcocb2V28sRof3LvyECfihiTtv1eXoiXS4j9tmITX2fEx+hJ2JENv
/Pg1iwKYpRqARRJ+YmUQtImf7cVupxrDUqiRXqrJ/kNETZrJ0hR+qDkD7GMspTs+XMuyodx4bvrx
FnQPiV0f34QTD3Z3kZVrJTKWb/3iSVIlIMoSqidLmhcts3eIOgPGm9YQvSk9tE44vQvwZ5HUUljm
Xv8XEU7iRS8hpoc58l84xRSt2voBVSbAUqNVausGewFrZBtJftSfnRO47/MWBVA8zQwxg0gbWuCy
RXFE8irBHuKsA7eWXhnLe3QLQUVXwAOaoWDkjPzQchs2DeE3iFzpgal10PZEoVDkTGl8dd22Gpnu
w7B9P1D0r583aMDPI6gRM81GkoWTjLNqd/74Pp4n8ou4OwenlliGcPw7z95CZTpSPl/vQ+Fk+4zV
lX/SRAaAXFpLScejBbpxzB6OQUcuzpyz5M/7P9pFSCPfBNaEoe8aKDjRB1rrYUsmSSIQknxBePSj
vNeSEcz/4zLS+FPyqgprUmDqUIIosESuocQpGeY4CQ6M6ju1TNGNV2906fJLqf00may+oKv271mY
3LkbQGqYorDXkNlC6pyb3wjeE9L2f6A/G29Ln0alCjTfm38/tcMeqpI979iYmH+NT8avIAHePsR5
o31LD182ErXZIWaeJQxzp00PsD0wktiAbk5zcA2xhozNHixTgc399LAF7EkX69Trwz2dym7H7d2y
8COP4m5WyWH0r4SdjDuOhEV940q1640ZvXa68iU39S1UZV6n6I9N8w+fWexuMq+PJ8zCt2ghcI5F
kWxFgTgiPAXnM9xZMDXSfodJJbSzt1Uj3ePNWu8mPCpqtPvzZOtjDImUUVAGZSPraoIqZtIEk7yi
lDnm4JvmwK6bpft66hGoQ3wfutKUmjXidExF5BaTttDkzGXyN8XAKkgTfj0JTVB5LOlu0p+OmB6+
iX9zfQ5njAiYp6FUAqhsMfcjh53X63L+JDoPiOWZK6tf5bFzbMyF4WxzCfifY9JHD7xQcKnCeyRy
t/40N77i8ku3KuXstqoCpyKYEPZj1KCv+NKttBgW8/PkEu8r3dEYemGC1eaCdAygP9h2oNyQolmj
+CTGXHD/EOkB2v/bJPkqLPsXPCkvkM+jps+mw81qTGwQOPc3lRnD+g9KbCazbZEMSemchZHKYDbj
4qPnfqWBIazCsJ99Hx4rk+NHXlTNmsousqEvv82ZNy4DLRfUxT2QbtYQk4iRLyT+xP1Jhm/SBuym
6QmCuRNGcsjyWIAM2whmVBy2tGas0JGorGyMEk2sdLQPDQ/5Wic/ZzsTKb9jCygKrz4Hg2r9cz4m
E+fVuhC2sKfF0BOpaF1FCuEuE1Th50fS5Gc0KswpZsK9nMKWRiMBrs+fcWuZxh7SxsPIuxDlE0kd
5Tao6NWDypVtDb4Dh19X4XnmN96BISmgWSzS8xHh3nEd4uZPJla9YKJ4cStpFX2n2LO6o+SDyMmA
iQW8UqIBVUk9ERkMyIVoNdnCYZocn+PAVMOLby219ZVlMc4VS51/IkX9Wgjv79UBpheLVkZ4P7J+
3SWHK4bgnnVv1Q8RXqc/+gSQlPg6aNaanFYUW4tK+DMIQTWIAxSw5d7n1iM8EpqsDjLyaUyQqJpM
JIby4CoBc4cQta35sZeQSP5RZIKZj6S9nAhbfKgh+IVSfi5dK3hQQG/XD0yZtL4i2oCwZ153pHm+
B+gMu3mk/dsYdFIV2tYSFSiCtkPY8PGEitQfJnP/KEItcLRJhFPVp/bj2U0ZKx7elTfsjc/Bh8tt
o7tUljarWq2iiQCQ0u3gs9M+Pc/UaTReR64erauVLsf/ByPRAHfRNWL2a0foV5fFBEDrxGSb2odP
xuYrAHFQ5a5ZqAxWrFRtYBte/+6BbRROJRZPN3rj5yjTSY7u6MSY7FS8lMbJoDHVhMwtMxcWI4km
2BDTditl95hCB+/9G8YK5Y2+Wzv5oj8M3i6Y6+cTOXO6EKZnGykD3VhkAennVc/ytHTMwKN4wmSF
Pjinxl+L4ZUFcgz0da4YBL3yQEh6ZIE9Wp0Ihj0DGt44giF1eA1WtAl6KMbBAaCrsHDT/OmFdXgJ
A2wb+cB653gJiceu3gALudDChHNTasG7fUV0ceGEc0MvWXUjzJkEGPBNdHg1o/5sgQ0BuUtPHFUu
RXxR/E3kucpaV7zYMCOKMKR8IZauvV9qheikllHGh1zTx6Uw4CR9cfAYvh7zm0w9TtyyBm6V0tKB
u8ZlG1PyiPiNTiGcM705n6qwiDdGYHehU6rbJB8+C+H4lhBUpnDvR9m1ypjT65eFgNGxWWMxfo5u
YQWS1mYY6MBF4ohcraWQXlzprODxu98r1OLAG3kjEigqpWpWddKokrJrWArYnSAPLcoivsuoD/SG
VnHpvQ1IG4HQ6hWgMXwkimoayNxxpM23V3H5Xlfttlmuw6g92n2NCvxeS/ABJzbV6kuWt60q+wos
b5jIwUL3hfV7TXd9ee8afQ5QiagnLHGwz9lHFbzjwMDXktg055rc2zLu51XlFlwtNtfejkOMu+gQ
TFPX3HmGeuqX7lbbmvuvRNYUhrKus5vfQifvsUwfyZbWN/NmvR6gawFA6RE2EvYFepXi+9u4RTIN
KctWmNOC7WfRVtGy/OG8w8g61tsGjVNAsPXf/DaLA3l9Bkx9ISOjY4jWiVAsyVilZK9oM0A/ppwU
s159p6TmlIDGu4RGKdy3hkNc8bS92lTdP6MHL2mevvOoetjGADLQZNa8ov2BRW/ymNexqOnucA2/
utTwIjmOOVksG3gaDY/daC3K/onMpyAo/ou5J0DCfYISMO4Cjho1tiVA5FbyqJizfL/Tq6NXvVov
BaBKVa3UIQxuB2uS9zcEvG5BVQpV/FLfcTd8U+mU71ZXTkrQsqtEJ6nZwbvmKiEGrOHOUWclSRfc
LqOoLN4Fppvt6EEfW52Y9kKdpBg44t2WsNrxd/L71lGSzRrjjYRznNgQShmpt5Wu7ixoLXXoW1Ad
mFIAA8gJQFq8zhF+HVBjjqLWFRFG28rDQ3xTBsX/L3w6/R0BBySXNdezN+ij9jmmQyJ68KYbl3zV
+yyjbv9sOFfZpMR9OufoOTbUC23atqvyg8Hc68wUksYkA/zWuqQ9qs+Ec/qe42m3VaCARnR1lIqG
pdzNAY49GJ4ACC3cUJ25AiL1tSthlbnrldGxckNrl0/DCY0In3ILkztCxFea+sQ4JaSYkmrcXh0B
LS/QPq7EK6ucjI8QLlJBPp89yes5KqJgV309uc6OtTdyvzmnKyz7UjdAK1RlsD8bHZFl2DX6NRi/
ONO7L+V9S6uQL1fyYOcdpt4c5ujfBgxd+8uffKF++HJlvg3neh0IVJLQGDGzFTk/F1NZuv6ulB7G
Y6UEEnPitFdY1jEDXfphwj8O7mkdIzXIfoLlVLcsadnNVx0SPZAHEvFBcjETXM1dfREhrGhSXSrv
v5rtRggFKOy76G+1WQZiiQqjRE30Xw+75zo0h31nirJ16wEYw5lAc24wcs4vfcJZHaqq/UGT4A70
d3H4k6EsNFUhYWY/iOUdNHYntYk+aB7GplGX58NypifnW+XTQ71unIjgq30NjVJkvpEKW6bskd0q
pCtzsvUpFL4QChE+WfKYz7YWn8GM+bFKdnRTxMG8iartDAwY7Qzdw81eL7jMBn2G7f8jDECq4sG7
5ki3+3dVDjxXasGpTevVSjioVxh4W9C6W8t7EqP/xXdiwshaCH6u8BFztEKPw/x/aSXjzMdJdnzo
2wSCZsxshfrzHZHiPJH6I36YsMmcWsxAQ+E5pqxGYuH1lNH0vBo/w3bsxPZD8XevcDJBNHHXzFRk
OYDtS1qUWdATnp9ZW7qBPjqs0sV9AmdvKUxivp+e2XJlZ35TInIUNSi1jtEDLxtcBwtznwjOHSiZ
A3ukWkm9ecWqRQfMF5Bmr5GqBBSYplwYsK+9BxwztbbEIpehCiOHCje40DyUh8jrTQy8i6lQ5f+6
SuLNsbfxjogzvDTMrcHw0BVosmpFfczjgL4EB38fBL1M8Pgt5aQwJnmZ4XxWGoGvtX19AAUifONq
Xh4IJLCpTzVAQOHiPPkjy7F6yWWVItRuZpwwv5tC45XHXDxxky5ffViw9fuVFOB/TStUkNLYiHqI
NlirqM/CnZvcBdmL+0rwzCv5PVOpQ0L2VsghU2rS6afhP3LiJTyN+0tfMv5iUlntH0DxmR3XLOz1
SyKrgWQ7KqLTm1om0bCDp4WaMpXEflW/e7U5Ntet5C/Xa++8wamOkpePKl2JD+g6gig70pPjCmd0
zmxoLWJASYiA8WCc/LYnoc0r029bg75C2shG27B1eOoXDOMgsd02J2n6IZxMsbRw4hfMlsK9NNgr
lrpiiuRFUSi94mb81fH91ofIXe7zVqzhqajyZ2sCOhIeOXjx3jFp3VQykyX/ze4ew9uzYBQc6PVM
IBOaqBaQQ8dCsvroip/GrYI8A2DI9zEX54MBfLKAum34R8Vstls1Qu9zNF7U6WHHb7WEMqWfeQzW
KZW+anuPUjA90C3heO5gbC2HteG2VQ57Nw2364gU4w5yYqwPphxJJehOPnttcoz1yt3YwR06QLvR
kAw569cqTPC3whaFrseIC5sZwArBQrv4GgYc6ufLI4iYFn190GclFmVCkIRoxgLQI9+4oSTMJlfr
SxE3EJ661tkQXd1rVpIfbG+h0VS9tE/8W7Xv7WJKwMDtefLUr3m4yXQdnMhDVNth8ovM0X+Mp6uV
tVP3dr4CgRg/mbuH5FIOmoxQAcSB3bXmtN0jC6ZEDVi4sNQenLS4ElgzVJNzOWo9ZVy5QuYQ9O6y
AczES9l5H8QXx9aYps9xZqJz/rprT7UkX77/ctw+SZQxaoShyDCrhIFV7b/exfJu+LLThiRPjoYR
Sf6sZfXb4AiPpaLNMdnRG4UlBVNoxmvzfMNef8Q8a11nHeWBtSXGx+SAtvYE50uqiXFNcS7No9Zd
TmPOvBzL3tVn923Qt5SUbUpzZBoCF+MLHfcpeXPYtkMjw/UXxStxBOIYiEckP+3bGjtneK7a0Ez0
p6zb22DrTltOTdA6uKcWOeWw7G2Q3AddzdVJQb+4TDUfwS1+YgTGugzxgaBVSrVtwYnZ/Os+/wX7
g7HXbUPc1p+XTqFNZB2W8EVJc8Xv8jq2jraBL57XIgGI2jh8J9p6kBTFl40MLkdna5FlNd5DDHqW
H+2SCOc5pGk/KU81V9YnKiQHABRNtPTEoQmEbOoG1LHBBFyIvZjPzZJmTzkwTH7VCwPzU1eniPJJ
OBSU4mmahcZfpmWnKnvpfb/COUCDkBSq+oF/FA9w3H2JDmuGvkJTK0cb22FYZtloEmvI6KbcWnQv
CrphfAhqBfpHRqv511kKyNfHXGFl5UZZtStAyI2Y9aJBQK7cHPR5IpihlzQuS+UkH7i5cnWNDLKW
pmzRdAH5MOc6Sz/eAwUd/bqpJRTAKPBPN6MtZsbI9O6EAM+tbJv72Yv9glyuIyhc5b+DAh+9HqXJ
q/bvDkPDmc9pW3d1MeUAD248TP5gFfvqB2ZpVcKHALvj6KkQj4v1C6rZIN2yZcWStfePBoBOLiZl
V7PA0sdfDp71T1F4B2ajsXfIZbbZbXoCw4ZWnhFGUIbGvHHMTu30u459vr24UiddqYBJ5Oy/08G9
VZ+RpDo7O4vPl3RpV+otqCWHBSPq+zjbZMJAp5/UlpV6Mb3mIAylWtBJNol0cIKqJ/Uke30jF9Lh
r9hPOfsD7/r5INyiJH6VxZn3WEdG4U2QE36jm0Qe9Fkwkabd9bGLZhUOl1mR0cVrYlT+ORcXE1R9
Q6gzUq7dQbTRfUIlKOZnai3aPuHYNvkZfdTGe0k40yNYO4U04IuCWBs6jm3zZRKVrhkr6587uWu4
IuGLLkA8XpafgBeycNjuRmQjGhnayflh8dUTrJFBZHcLnXPalUl6IZjDgPbYekXFoLNewFTulA7j
dsruDBhgHVzRuNMk8FdHST0Rvj7kqaOTD/m6PbzsC4cXeN747xJBKy+//GJtUak4p1f3IyCIxlGP
roy1RzwiTm85rU9p7x7RBH2QPbM75OUF3jEwb12VYMSXrLymBf/ah21mHTOFaaRfT11RR+TEfjzg
RKhaLNhpZr8bxh+1yBkGS9PvRRu7qYv5t71N2ZMvlsn4iPjdb4qVszcRyh1uUVgWOB94/fOyNtXl
1bSsevtQRjQ8KKjKxZUVo7e3TrYnMI+6FcvSfZJRR9e+5lm5aGMhgJ9/8c3uwWxKIXGpMp1li6jc
Hdh6rhVxP0UqCM5vnW/J6/i4SDES0hWhTSH1dd+q/KZCF5zE/E0axwfLKnsGTWXNI3pRPYoHWuAi
/DH86Xt59dCIRox1WrEN96LmOneFuvP6eqCXC+id5Wamlu8aezzwbaNXtDypxHcRSDWXK8aTnlmv
H4VouH1Mrv5QpD/JVGAraHkQIhiStQi1E7LkMB8gM5cMZoy9+m6nWMNcxz0039DXktr9eIIthL/A
gL52buzu8sMlHCj+8mnxvVF1Z9uFS//I2fihhqAqRBAiZ1AFFH9rx3zyX/DL+hgDCB5qOBLiQ0aD
M+12hIzBSpDuJMB2ZWdTN5u1kKDTqjpEvYNh18bBLp0h+/X30ieSOQjB/oVKfjdJTOqphGDfeDJC
+hoT05rbmUlhW2PGUhmKhk0qU7U5syir84P0WvK5hdQJxyRow9bbFEP8YxqnaGJsZqS1uKgC3atv
0cffARQqAraPLAD5IU8hImtJu9Zfmc+IDdmYXL6Fq0CNo51CtVcmFVPOT59JlLmr6wHDL0xx68xX
zhu+TxB89D45JCC0cmYoSLPM9HOSHrvg5/rgS02PZBuA2XKigY7DBRzE9Z+ZnR/7sXwCI8t1mzla
Pty1RqCPfenAMf2ME8P9G+pfcpq1c0zRz7prErHzVel3tMb/iMH6aLAe+f5XjaCQ4jpBLtA0wOMZ
5idClawdAx4tRND8zPT0qOYMQ93ICGpeI75OCDwXVEDNekk45GN0SUXbAnnrrAnqlbbNyjsbx/9L
nugWPXXnVGTMXy6y83tfA0ZlA64vkAd1Jydc9M99f5fupgr0gmua/t6D1atG8Oay17cCE65zYbII
KvjloVvtsjS7lc2tum1Ba+5p8/h4NtLrUCo5zTuT4yP42I7o/Pyxx6TXdHm2afj41eb0Hm7t3h+t
zVH0HBbhuhIpNMJUaO/z5yi6NIK+0zK9R5nsPul8h6ndKY2fBiun+rdowBKoCK1nMa7Cu9+A6Sjl
/QnFjxDv1FIloTpfVB94MCRjSIJGv/tuQJ+zjpajaCZ80rvyjx1Nnlw58j2Sr8x9YJxxRsowYpcV
EXJUWvWVivZGA7QVFWaUg2hhFALJGvJ55XcPWv/1DSrB4+z4OxM/B9Eiws9GYz6CUlgisMfPd5r2
qBg42Bo0JFEiReSwpY/GlpbdJc9uDY7VoiumsOQfqC99f4jppd87cKrjuH/n2jDValO69qUeKl1A
3g9cEG9uvzA9dAgjbqLaWa3crkJ+kBvmcG51ZenUF8OfS+PwUBRsv97VPbWbldk0Yfyf38yv5XjM
zWKRMVZmbMTRfa59h0ztLOJuJQEgC2rnKQBHhRmpnI4ubGaU22kQrI1sian+dVaIRepCO6aQskbz
VQtsxLHlaRXli4Hf3cc6eF1tTdoPsl6tIBNeuDC/LPlfThValArEaHrUVOOGk6feOLZMjTc9aaW/
U56PMPqGtXokHUBh6nxLuRgmVUSt48OjQ237f2756Pgd3ZJvW7rQL3dLlxmiuBcujUpmOAMOcFka
Sz6oJ+2Z862zgIGvE8KX8mPlHYQNs0BDtu54z18CrDWC+XMf10DRIMwqm1itQLEyGp5P0hRC8QCC
r7qp3Pgn+WGrYxVRphielqyxjtZvZTlaWmYslK4lCOgfDIsrlfb8oc0mpyNV1kIEpkeaMs2KevU0
F/a2ppzEjRCwMxE2ovnYe75KXPUnWfeCCvEpdkCQentJC0yCU9uByxXnto9Pe4lOGS/1goCUKJ3d
kpJLF2HdRkVUPfc7ZVbXBXrRx6LHO1CrP67PKGCcLh1qKp8AInONmTnw89vdUAF38hsqMYEueRUp
VzUOp6MtygBVIqEHAA9OL7ld1X0lQ+qwTWIQBHk2YSuIUa6JdX91F9UEvINYvXZFBMMsCmfTRUl0
dsUfTfds9Mj2T1yOcZF414ps68PvY8BYesGejPbH3MGk4K8shGBwylPzJBNr1Ons4f44liN9Kld6
8tZsAxw/ZBFzjU/P2l/HOZM1DteudsmLOJkXwUS5AsUQO8xcL4NP8TMdvTkkzYTSmNNZFMatKh3O
9I6C0ZoOALFibldi/5T5JEVHRkbN8QSAjlmI22X+DO7/neQMMBhs8Q6kaApb5oWSvXmz1zUDlTr9
23cB/vWydvfs/gMkAhNbYHP5HgoRMcT9GLEIOD4LtsuUwzsoy9UCVCmXn/Ebz3a5kbZF7bxsQ9Yh
aDZDkL+6lfg0XBmYhFjx4ScigF9nCuMHIOJZ5KlFRhSLtJDzy6N7kBXZ3CPQiN5V9547z33FQNJ6
ajHwqpqKyCXZHil5S8kueYNOYUH6iN0kHbbQR/3dGJ36/isI+Bf+DPyfieNth3lHTJd+5cPY+2j1
TPHvTbbIVDA0qdVZsV8vmu1GjL6Wl7m4m+nLxf5bOhO7Urnq3/rSdpryW+f6zn1alKO6wBt8f738
sLrRwYJiIGADg8T9idz6Vw0mN5nqWLTPRalXbC9oviKu1Jrqgj5Y+qGTQq5k3Eqq0QrPV4+AbijQ
1JrWoz5Z1lulKl25SQhEYpOQAqZ03vpGGlFuZO3Z7YlQTSN5+blghQ68k7z1hYLgB2J7lho/b47U
RIvVFHAO50jxGxNzpBaMVg70fYnrEi7y2p2kXOslb+TN9yiQeai5iQEqsItZiDWwp4B3+OwG2imL
WResHHQKsiaPDjUVKVGrZsjEohQ0Vb7WewhFAcT1n8tBLwyzKHKfTnrc3V9gKHrY0xmmWLmWNmXZ
bvey7AA2oKqkqnNkMw4Rcf+9IXuGmmMF5FUia8hxIfxgo1rYBwc/kHGtjtbyX3IFoNeVxCqubpBs
uNh5GutzWyQ7hFv8miNpDDp7VBgY9+zFH2HDSZ4Ie2usdoktJIZNgLQxU7WRvpmYd58J9GXU/9wO
BzfrLeFlDJBYpZaijeyxwP/jNTUSAsIvODaunSu6N5Y8RfwcMVRX5YDyGfYDPJD2/9ChrkKwAQhn
zskN63zDUaSuBvsaavTd/8zAm80V9vS+FmziUodOMFx45P6UfEaghNMKE6PA4iEg2yKgzFJjQxTk
t2+Mz5/WA2SWNrVKQ5kvPHGKs1F73WvLJU6FehkNVTVJkdkPM1ZlstSC6Dct5W7xwBnln+eO9JPQ
GEtvannVuHQF8YqR9H1U/T/mO3w7rBeIVIYBE83hWM20IPF+GEP3ZqQYMg8s5hoyvg08DvEkDOvW
wrVrOAX8mVoT9BLhmVl9B5UuWVgwQilt1+SFXLdHNWczbLaprZiFuYVecivIHqAaWuaWa9yjpR0d
dIRDffGgJDSMWLMSTY1Zl3hkqhNAw4JlNMrRqHm76gITJiiysIhRbJ5Ib6xHjCGF0a4xo8anNExq
8Zz9rQy49Cypi/2JaJ+Iz5x0PuTFd6M9jUZZPuIWJyQ/xD/cwisFivz7IqTR/W7QZ43cqxZ+NEe8
CtWK77IUigQGf5AEcrLWUc7dB1A0Gd1oPU/9obktyQL4QRYM0Eta/qeMQiZQTZWyOW9UDW3TGyrD
aDwWG0/y2m5FRogLLdeVLUrp12xJjbxAtxH3fL1hrj8dHeM4vWLIyyL2OSigXNmsxWA9JxTeHB2o
en+C6B71eORZNcr0BDV420fL0xmeKAPxLM9DYFg5j6sQi4hPEaDusjAx6HpoG+Scn8JdIrQBY9M2
pXIzX2J/Xd6x38Cn9y32qMgA8vuf231BaOEKd4MjoeMLSCha19Y14kzOgyvZs1BKEM+KstO9TL/9
dcoDYdOhjRkYZdOg/YVMUuasACAVj6mMXnY1xoajRlrrKCIZ4xfFyw5jhPwZiKPnZwe4S6ZCTK1M
7zyDcK54T09kJKvANwfW/yIrKT6isDCS8Yn9Wk93DSppFi1XEXuXWyJm0oxaIMIPFstbncK+XBsZ
oMwy88xrH//t9PTzNkR0KbIi203gbBoIQIuPcjrp4E2nq8uXbtbkFL6ZxeaFYqtaZvLtIlkrUjer
smLfCMKVOf57SoPa8T+audT48rL30+LJkZjguuplsA6OrVKxc/83L9+a131gHw442TY9rpWPpQ6/
Re8D2vdBsju72SzcCNB0kjhBcg7A4w1r0A1NdsEpFc7setcO2ODpmpHYQSu0l/c9/kF0MSkTKZ73
qZ+Igki/sNxx2dWWBymFeUgEa7yWATVjh8bl759g/Q2WTDIosLrY5HMAJspLSGU1zSrGR77Sc0u9
pPWFyoQQ/u3LIc9GvFkXia2nwKwAmRdhEqQIW5yRbdUjLQqBJudRvJUKPvB339zXgQBvu+Ezu+Ec
HZp58iosth8xJRdhqKs7YSZh0MSmz0jK7GwKKt1z2/UE7tMCpIvhPYXAwc1lCHu6DXUVJ2HDHFei
6S8SNQHyW8HzHwZ7Hfhaw50tmCJmPmZ4ynQkdYhn5bnMoIgsRKbH36+cDTwiuShWhEv8IXMXUO+e
dL61sHDMpjfeTzj3HfTkcwSZrv86AXMzqHUKKB1O1Arhpt6bfcI4AZOuEJsVIjmQRM4taSNZv7Po
nIKBOV5RDsPKR56thvzlsJvPHKbkQx03RJ8wsnAYkbdscvUvbCSMYlBJRtI7452lSzPTnrmOk0FH
K0EzVxUTquqnNX7Fy3ZdJQnU7mZW5Yv4FeBy7ldYMOsWyDH/8FfRTvCFEhXxjybtdblrTYv+7Cp2
KmurHyKNJVb6o+kHWBBAbCwW+pPK/pM1OgWrMdCwxxsq1WnICR++VN/g63QK+AFBMdShTG6/zhm7
ki6iVLhHyD7j5GRnODeNvrarP900oP7wBKUDbPSBQMYF85lzyXpZx8w3pcxkMFozkjD3k2uFEqLh
5Z7wN+Yvjva2QNuLRcxiLXAOQ9VuhRDS1SJt2hdCdXGK2WvxTVrWD1M0uOn/DDwbM5yXJP68N5Oi
gOKsHVA7d5EfO3wh9F/D2yNDZYpuDDOJG2T3yDrX6/Wwj9dNOX45l6R5+uP2Lo7kzIfzz9wnU6Wv
zjdlS5FHueoqkhZlnj0pBpvaBtQeWCpdj/RpwqUE5O0KH2d0xIFVI0kWufNl1QE6e+Gqq0RxULpt
xzDFxkQXLeWF2dXWbihel9Sxdq3JHKG+C1wlmeXXb0oPawBX4lFRjfklPnwv2Miu+cyrxIV0tSHm
RwAU6GddjdNqYlU71KHe/CoKzLyNzPAEAFFQ0OEnQId4YlOkSEOnHB3VYX0NTT437XIk4BZZQbhl
tqfkPlODojw7hkQXI6nSPplsnOWSZe6NPkyNDoJWVDxv/141XUHwJkLRHr2iKTY/ukWVfEQpGsy/
/2kFRWwBZFMPHSbyxiOD0MatzimT5dNPuNIoBjt3Zavq4XFXusAoD085vwl5ohTc3h53vyfhGJbx
NiwvIu53mxwoe59qgozNuZMgGM/7hrvE5vmuKa9hDyghsN/6r7ITjmqYbQV7TYzCdcsmaq9mNSAf
0jrWn3v9Cv7LNfmRNlc+OGyR1wekv7j+OL4c9oyNjXaDAH7HF1c9cLaBbsWzj5Oqt+XxmFCCcq8N
p16nlVwWRcx92JY+67nNJnbqbmkm3iNVRz/VKwCrBQ7UGEFbCm8vC2hBaLPAkSYXJ2Qj7Il3mdUU
V65uvTcnToSRfnGBKYmu2yBveTIAjYjficOxXE2jMT7/Gpp3NN+QdEZfr4+SZw1AIJuFR7sid0MD
BtD8DiQsGj3sHs1Qa7OcFsJ01P7KCxHUg68lWdYr1NZwvu7ylAh4lfdY9b6sQuia01SnHAtJpi+o
L/tThSY0wer3dXTHE43HsK3n1VT5o+JDtcF1/Yllr4pR+seDxqJTSsV66YPKTk4DlC3Ut/VuZGaF
EshtvjfdLOy13PDNEPkFIo30K8MrxHL8TKEUS2mW96BdpuC1xClaVS1rIHpCtZcHGkmObmN5HGrF
uheQCUfz1lZSjeSNKnxiLMJHM239101JAbdfSOVzQakbiJ9gTtZgaaz6AaNKmXWXp3D/RvIW6xvr
1XbABn4OYlfVPW+dzOxUoN8n1KaT05ZwD8AiAawE7bh67DrNAj8lz1hZ3OT5FGRWRy97hUuvDXfa
XQ3LJgkHj7fyzkAJAGAfs+fdf5VmNU2TF31qTRB5RTA7h948TMtOnrm4HtMQwkRCrNyCVR07SZQf
G0r2uHB2IXxQ/gUB+VBRez20/bt3hCx+ofe145OXi6xDesysSRhY24rpuuHV1Vkfez8zrOuY5fu0
nswZVqtuU8GaTB0ziTyYoGVyocK2nECBkkVo4PA26JBz4CThb3ujEJ6q5+kuwLPfbDFsjBejmn7W
jps6mWrqRcB0q/Jhr97Gvx8SaT/tnW5Yjh+Uj+uRBcuYvUNfd63E3yCPNbkKRtaXceZNxgdrQ2Wy
TSqa17ArqqBDn0d4+kBhDTeL89HPTJ7XZL77+01fCRor9GVcXi5+/iQPB8vs+RYiP4t7tAPV6WCB
CFbmlOIQiJYPkXYRb+8ff9W7JsARGEP2wkNzmhSo6LlH93YI53nRLKTqwrD6ZFL9Dj9yavhfFJcD
TjhZdGQVy3RFDz2mQNVc2jmQATmLjs4IFhPb8DNIJZ5qgJcGlFIF26DnrCNbKY7IMl8Rxr3ax9Hq
6EjXWk6L0HIDau6/N6S7BAxfiowSy23IOm5fhEHrORcC4XQqwNdA8TgGYM6nlDkPETI44x+vXDtu
Lrei95ti9Nj+efRr5g9UjVTTzkD00MD9X3Xt0VsZNDxC23yb41nWjFw0WbJQkn5K0ZBA5vKK86W5
Fg0ZzDBv5/f6m7ch1d524lclr0yLYKN3g1ccSP8W2Dr5QdVTGHH/hjwQvc+hLg3KP0x85MONLDqD
iS2r6BtpIXsJBjZn3hQI1+vpRb+2+g4Sl7/y8fMGfc8RbEKltZgiRZeLMTMhxvONuGwtQHIo9y5h
XQKJo7Gl6saXtRMMGNNY//G/ESJ0YxlX8y2MaYaF0fjX7hECy5XZ3UAFGhzuhecXUC+iqPCI7fgU
PVwG1pJX63Wt6VRNpGHp+PtwyvggwrFXh/Am7PGurOYw50WNiHj0jfREgzSAPWyXXs9SO+2dVP4A
P/gmLZrFsW28rrjZo45X+ezrEwoaLE2HXp2o5WBjarWqJUg5vOyOXZntXga1RKNxrSBmUYJkVNsO
5PMWjKZENYxlrhEYBsiDRtSuBJEJ51DkDgI61eJfSzVp5nq6CNqXdWusGJ8mrtCP3NDXnwo/7NOA
YOH7jbuwFgZHdqpzP5ZJyJa+pKAZCgph2394LuklrrY6DsTnB2gudEybcE6ATndzUwbDx+jXUdTY
GI5+M5ZEvydoUIPWTYA4ir7FWUXoa4KZCNlIZivhKfKrom7Zpp9ng5kLrvWfHFvqEUpO5zYKDZ6z
KMAmg1+ecXOrhBYDnPteePRPqeH65bqh7bd5SYYoxlgPfueJleOc4b6GsSJquEQQ7mFBgp/CesMx
c5ynU2MEi32Bc9B0L7Y0fSp29yVBgnBnYbbKTToo/cSXXEgG9vySmVQuMVVa02/n0NtIgGInufde
OJmmmZc1A6R/0doQ9QIs18RSD4S1E1Q2wciRCL9xEVXD6dXUslbDI7fR64nNskZ7J4PLvd9eDJJ5
uffL4s/bJR9l1Y9fejF5H7Iky/y9/UkbUFEFVzW/pYHaYg0qPyx8/nNPwh9AX5r/+sg4NjIaTBG+
RFizWSWIDsUFZxSJJBe+T3vLHnsk8mlwUk9KHGAEK0M+3T1AEE/r794Pia8Dbt2z0llAccDyq1qo
OcYsI2aAhY8L6WPnCt8Z8v6gF/dJKH0pECGZYzOKiG9XI00FU4v0MstmNDLGGRT9n+5tvJ0fdxRz
6fVSpnZsgBocZG1JClnaFAxf5z2on48aXluOhA7xd/GUGSz5kA3/fwNtTmNxd0Wqk+ECcOtdh43L
P30iAyFMyq4xDVmqVGu9M+k8YtjTXEwc5mr/2KIWxazCJ4pCt9lLnweSP1nvAMZwRR+r24MRuVto
0lVEpcsmGfLdxKv89Ec6n/MRi25x/OB/8WVBLZgt4DKFWPBEsXkyFI8dfvbVz3BLVMn43+62pj0W
I4BKCJDXiBhHc5s1c4Nk+frn4kEzTNNsGawOQ88bS4PRuVS5Im4GX/GPpLnsXgvJLT33lo5sIMa+
/yviugbOW7/8yHWVDs/15LOOhbz7TOhNXecqe2ip1oP86Oh05+rsCDGwyuKCAi/Kw/pL9uXNOR6x
SNi712es9XBN328J/yvmXRte6cxP6+dNKvFjyaxyIs/oDpndoJbsNf8sGiXgFzYUjhFcOKW+hEVN
5Ryp6pfMx7PIWOZsFq0BMego8td+cigPXx2PWU2gFwJLugKYF+uwEc4JgDxRJ+0Wtjej+CXjL9Qd
aoxxBfIgzCdI0REoX2AlMZudIvxaO0C0G10QhaYKLZAT+TIi/jX78G1CTnckg5fhXwAp1YrjUk9g
lh8VxAZRLaK2hnMmFS6QGAMxAcoCzip4LYfitjKWZ7DK/yqIIlp5Hw/QtCNzjgMyOT2eRhKe4C/u
I1sQdwAbjtXKR9o0MxjqFitLNnGzBTmizlpzbHoDOq8uVXqZ4XDUaQm3KOIed5clwCIrDI/28ZBG
vyUVheYC2poxHA5JR6l+bmIXHM/bKbaz/dw5L8JnO5R7gufb9HuwiJtmzoMryHCWA5UJx5Uet2zK
1E4UFmCvRvsu3saaRcClT2Pq3AJ96xhstFq20QEWojjUWpBix9MOY/d9injeZVnt4hgGIXTCYBJ/
e424QJorWODej1MDAmH+ybq1fKP6FS/ib88AnlJA77UhItEmauIFOkpbTBZOGsHJ6DucIx3Vc6bV
W8IH992ns93WP4fNK/ZRoGhf5hWnMFMnoyeCmJpO1gZlH9Rikg6Ftyhe0Nuadk1YsxSCHl641HG0
wIMG4HBIVhIWp3Cmw68csaCmrwrrhUL3IFsVIWF1D9x3qYPahTymMmmFLgythMdLVZwjEEKGPhq9
uatlxa3NvVsvPm6JMZNd/V+TpqrrTzMR99fB/zF2KCaeQyue0BlzjJU7puxs7G8+5nWptH5pB8aI
/4MTnnWKpCae3Qn6NnI5VCXWmJlsJqe1608Bf1Y0tyoT99oPDWWZI51zkygCoAC8CK4jz1xg8FXH
T/H3GVStdcYKgrp1bmb9UXPFJ8wuqb0xlS22l9gcgZa03ZydmJfjjrh2zhP8V1epqEWzwrXkmS70
Atl6XV+AO/+vVL1ms1nY9fc6SXbssLX6Z5g2oeP889SGtm/LUQ8+JizevHXCpimOHHi+CPt4k3+Q
GS3ch4Y7AmbVswhwSBuFTta4Z5UQGumXbQWe0QyYkgxcz/Xcw/DjT/pUcMkbFxE33lSs4xdMCGep
9Nm1h6/11eYcf8XQk1KUS5sSB/HK9+aGYyU7MFRpzfM6fVG1Mm/FOLJ/QnVfnIQvZXq8i2ImDNKs
GEG4L+/WveCI3Rahxr/if5qPKwiJZd8/q4JtZokxoWmG4FASFKlMJ6PYihDRYO+1gNXgb+719Ysz
/d9aXYNENmCkohemCWiMPP9fGh7T5Lg9gc7RSKsIHcBgOWV5zjwZu93lr1vJ49L1h2ZML4jAEmba
XehIPxuuO8NH14bamvjKHFo+HFppN4zU82w92rrtTkCZNToDrsindBBbrCPphD6LpiMDqcWqQXdk
WRqQSL5CoZhs+D7gz3IyBkUtlzYGokdYXWvSIAKxtdE8lsvnOSereXKqFz0IePugC3jINXNPX+rW
C7Hek+e6VlPz6P7BOY2ZU73toXiEGFcmw6CY+A0VYZGZ1QdC4W3ERuUgB3l4nOxay3C7K0GIW0Zg
PNwq10c5178kVps7a4kNWcMlv9pWYvgSU7zpkFb0wKRv7oZYIjp4Iv7RIL2IaQdtYxvqK9PDSppn
4T09H6nTAVuKU9jcINQJ/iIq/oFAREFHHUN9rKtRAuoFgyq5epI6nQVn0lcQwYMHCRTGb487JKyA
OJMk/5vpa/yMeOoXbbnane9Yj+MQSuGusqvWK74ywWLdtiIFa+6FZ7l9zBiVRDAhazjNUZxocyPB
yRrgl1j+xeJol9uhoSctZIO7F1B1K0tL+5kCuRCpISJRy3dFhniPY2I4LSBEHCMRUdBgco+QPOGW
Ps1VZvNT89Pd9fJ8CIpQyDMOHziK3p5Mtgh0tmx3JjqmFnfvtnZwKNVsNmRDzjpqXsNoWd2SFYUM
0BU6upHYYF6ExB3jxGZ3whRT9uhaaRhpB28rPvE6i4zfGphwWGiRjslGd/S+eqM392RepP3Iy7cA
YpVP8qMFG2laL1jtMQLMIt0TGDF/3BQWslxs6iqSjGAJSU+LRq8XeT7F85G3qcO2giDlb42rDcJY
xPjcKH+yZJhD9Y/k4tpmoyk67OZOlRR6z3jHvfIy8yezC4QcAQNDG8V6/cNEl1QjI09aEIo3p95N
POmHICdLcPJ6wQfbhQWsfB7ZIUfQVdDYMy/WGM42zFFscgRe+N+iCAxmjSk0SnDpfsRGPIjB/n3J
b+bp3flEb2PozLn4w0SL4Okl+PLZcR2V2pVI/6kAkJAQ36HSMNb8t0KJMrb6E7t436r49tUQ7Vtu
VWhhe/7sVaSdmiJx35Q9huHPIQh0O8NauuMSQAVyQUyZNNCcN+aoYoPqP8vuSs2Ty1zBs3YLcLfH
xsQpG7eqbF2hCNABUIG2VjCyHsFeywOmOkKrZcqwf7vlrny9wlplTaN3/2ZpOez1UrOI+uRubn4M
Jw8bKnbUsZ0kzM/Ui8ptMuKNsIKmbEr2R4DRVFx89Nuwd5INkeNf17z6oQe56/Az28+JQZo8Q7m9
O2w1yqO3Q1P/m7DePGhV4myRT12QHaFgPGa0WC1eVr597qqc83h7LB9mTXwd+hbLhy/L+K9Kbp1C
ukdDWGdmFQ7BpRwnrCsfPK6LvqT3gtDGXRsifzrpCno4IpJdDdpsBymQybdGPxE3DHkSngUHr62w
FvVagLAiF5GC3FQ/9z//RAvNm//Rf3hqYPGKUe8XGEtlWp+AN3SHTkxtQFBZI8ycrS0JG9KNSWug
dvoiHTwtgFfUr19pSaKwCqRaz+gErXlnGl+NjDO87CJxanrL+qVKhXXqy31vnpBvn+C0m4sU1sJh
mOK/NFUutt8+Xnz3nDkgAqbXTt7I/P2ozo5LIauNh8FjG6M2Fs7ht1Yam/y+fUZAxtTCS0BimKKY
xfRRkjb8a9gJbs6KDqJzxd8cx6z/qfzKpWrze5WYfGPG9YVeiXbyjT7P78fX6Jo1coSI94rfAeyH
KwNCViT76geXKqKBZVM0WpQe+waGptaekehiaB1itFmvI52pvlL8w/CXv+f5ANXrss6X+p0NwCW6
kIvwx1wCVzJMuVI7c+pM1bisxvtIls3Qg/20LlXxRiaQ8d4QCGkzo6xEU3ArcuxrBjXcu2d758cz
iKn6OdjIVrm8xm4Por41BHYO3+ltAZw2tIv0T7oCLj3zyVfynZdoPwZWjWfBoWr9DRqerFkDBU2d
tGzVEAGPUCnpb2era+eIGgLf2sIZ1DXzM948SR7g80nfodfqBeEgv0Fk0TOaTZZNk4J4lST158hO
p9EIwgjhtNAoiQKjNRctivUIffHRnBwDCnIkzqtJI0fT7mBsx7VBuLNStVeNh/xobcoc41mJ94P7
RmzZ4u0D+MBPohcbbfY6f+cdk2MBOevDmAiy0qaNq8RlV21PLrNbu49tzG9FZStPdOpwPtDSXsgN
itWl2PuIor20e2vZRxq5titIqOq01AADH22Wq35D8AnCWNJwf75zObTLJ24UaspaQYvG9h1FT5Ug
w7/9agfTQ9a3iZDECDUXgYRa4KJC3oczo1OqiziBQYD5V2EqL3s7bHHtzaRMUdOyjV9EPeCkKiu0
3mXPupFQfb/ZuP/8bte2bURzVaqPmvl5oY6HM+2/2xdQp9Np14Esr4lvcmRihFUsVScr8htP0sCV
QWIRSFlHP9lYBcd+P0dcb0yySw0IUB1ZnWu2hPb0PPjJCP9khxkUQypJS6tfBQzdf1eGtlIwmVHh
hpUcH8Sy220vyFz7ooRR+RaARelNnEusynQcJzA2sWwj2EJxMyeh3hd+b00vCw5KM12pGbT5eOpG
2u4WPADWqRyOTazqK9g/JuqWJGHUiaiYvejPsvQhniNwavsUddQDqClHWVgMPdxmx1+ZEdJW4Gc8
mIbTZrpN8cwmo6hdxn/+jIPrKga3txWh6Eo1GGQ7vbdgYnDPKkt5c3ffSATwteR1qD7LkVMEmVL9
ch1gA+4jA8+ynR83js2OKQk/gaVvWSDgByYJxM4HbBxZsoG9PfZT2lG8kYOYqrJJEfi0uUNEMGip
1tREZSWX3QKDbO8nigX6WPc3PZ/uBr3TOTwO5CZk9hwKkaUocIPl91MKn0tpdrnMjOZPaY7+R2fj
gIcIXeKtO4HoinPzIctl0K98WTzzhZufU5fHR3ipCE6s2AA/w4gFKWf9ITyeS2z+OmCkm2H6PkIt
EyiSPYNIsXaP+pQqSrFbFATJhBdbePqToeq1DImVyVTluiSwJpMS3V6spZHZv+PykoefHUEO6O8u
/u3jjcSsb4ecFuueMiObKr5XDWPL+gI2CgkijVgVBISOrsG0KPoGi3LDnYO16lWndHTI1DldMJdc
CJb80+krDS06L7jvRtwiQ6vX2CQ5vPFYytRvgD+ZZIFITFPdqoRaTUeP1PpECeU9nm3d4EIh8luW
7PtYg1niqgiq0R4RTRPNpCTLo3HcPSGN59SYr3UlCr2i2LQb3XuhNh2v2leJ+hHPgHd8CBtSLWH0
AothnT5UWQ74DlT2P7HyJ6sftMP4fV7bCjt1GqXkzLPdeveJXNIpIq4vY8OLFhLrBiQY33ZAVjRd
XUHRuu0kNDWgTAeP7CJ9lQxWRDE89XTQEDFqZxZ2m+wxzSxa65+pvbGSHKdjnCOpVM2DtcUEOZO2
uaBfJTAR2ZWGPxVO73LfZWap2diIPsmlbG0tlHYMcTpLozwHXf39bX+SLobRi1/bOh0WIs3WN0bb
8PqZ8wNicgkT/2hQE95KugpMFt9RQIAuQpRSMwJHLs8OTPGIxho5kwQmH641blrh1OsLtXe4SYOy
4vuDlGvCVNmABMSKfHkd1PDOo+RABW1BTaU0yn8CkFXYfotDLyWMewmAsm7qRmF7zKKNhQZ09nvU
CcL5lmPkiGGcJhgpwlW1XVEogSFIXScR0B3SgIWk2jYfAm95YluSyDrFOZXNyaj3AtahWbs7vNS1
RhjcMEBH+Gu2bDwDJTi1I+Lj+BZoXf/qu/UuXL3SdjBWW9SymzZIeZ4gXpM+JLeevUn+l8Bc+BM1
CyOg2FR96V9vuuSGjJLW43OXg0OXX5sB9txIaR+Vo+A1Lw+FgQQLkHDkiG0UQ3tHfdjQvobY0usr
0FvBmj2jg2iwvRQUSrUz1D/b/0xYxqSeIpVd8LZRfNTExRVLoLobX6p7Phaj+/omjnKzhLfT2Lal
HPMopzuF7aOk3RVlr6ugeAcUxa7LKbEHZ8spOpD0fcz5B5/hsYVUz8rjlCIVO/5nEXXRuO8g7EH5
3YoS3/cBbQ3WrPJ4AzMSbNLXCQyhdRsrFn/PPJlhYCVm+yxvOQZOs3LSr6X5D48fDr7zlx7SItId
BUABohLFnpohdIhjrkGESc54OWf5P1K5T0ZvH0j0FaNOFxNYD2/wxugo/M+up35jWL4a0DK133oP
ys2bWqzUU5IFdGPT3r9EUAIuXaMkWvtapVbOsZuA89074FVn4kRFc+AfjtXsOpbAgYg3IrpzJIMv
4FuLO2sYYylfhnj7O8lW1IR0J83pC5ulqZyFEcwXOXOHgnT6MorK+VGq8b67DHHWY401PWlObw5s
//cdYuaVEOzhyZoO000C9UGraGIz5qm3aptMrnrX6g6I7knTWB10XXbRf9M67q7VYp4xFuvhOe41
Kb2mw+IT1mbBNKtdZ8MbEn630hQ+2IvfdSOvfCqQFNt2kqkWofPhRBZQBexWNw4Bio5PlZm9YGfV
dxP++Jk/RM/a62quFqZ6syOuc+6aeob0Pse3x6JD3oSMc7KCKuXAyj3V0/KJwdYVE0UjibbZ70LK
LrjUYUYHDsr7SabME/o/ZjIZ90nbYr5pqyaD/2sKqjMDBFEMitTY4xqfeQpzIva7dfS+EvopWwjB
mNvKhpNiANe5nVNjc7CzhiiCVgu96s1Rmr2hy7GxGdLHu2Xsi0cp4FwF8nOlOkZCpGjnXRjworUk
cCV09/qa84DVGapAs59L9gJq5q1RGHayMNhR7eF4HRgn0tZn3Hl0I/J8gfYlASeJ+MiAPCI1qzkj
rvywKwluhHGC4f9+8OO73OpYoGvH1FAwpp6TmFSsEqXjX76DbKOvurgNUoj88zgPiBKrhjH9Zfji
AE9e5LDCXf7jxyhcazHdfFMV1VEn7hA8yUQrXm8vK89doSOLW8bkqhcX0UQBwR3W7JS9lZCwd4zJ
FTKRx8sqBu4oBOxfSmcs+IlF8xbYbXNWrAqMLJjy5W2iyxyogud4qRp35FbQlk57+PAYgqOuuF6x
HBeyKOpz6oePp/QIr0XEFz9xaDEDpvAEbgrCBi3tJ/KgaLfGHOSKU4Cd2qFzP6zJ8ekn/0mcTZth
wlFyM20urDRJmWU81Pnew9CseZMdQBCBfosgwKrPxGDEficUs0VejMFjA6b7D45Enk3rVjFyI1A0
CLSM92ErjphQBIEJXcIMFleAGeJQehVhL1IQ0569180Y0/TsXY31RCQCAcCnZEELDZW9dGg4i9T2
vnSOYtnkfdxOGHkF4n+yPBozTC2y76gu+FKOkmn6ICHbwrScLk3o9jW8yrrhxdEs7/zhyNQmvR++
+MvA63pb8FeoJfN9L3TrYH45tU8BOIvCfJu+WfJ2Mf4mjed1AMGQrSiCvV6UN9ySx4t5MegNpXKP
4/qujwEMYHdP2M18v48vE/6FOP7N9IS7GEq09JRb0+3MW1OFglF3FnRIHEFI8gbTj5sBOIXP4/UM
NlBD9jNYPIZavGj6g8TVb8ws9WAy/mcXCUzIwskACdmVpqbItifUZwzYPoQ3ByzdyqsrCQV+87c+
cqMgODk3g0UyU5QouH3B5O5bvk9UGqGA3F7CwLhdnSS8WqhFbQFDxpkyZFIQBgjyn0sfwgq+HS4r
bxPlva7te9jHCTwMERXQcUPqAvPfmQFh+hGQxp4+k9cRDOKLvjNVz/qPs96PLu7jCyrx4qOf3j45
Rb74Jzah+afG3gu2YPWe9mWswl83VhAtS/qUpkEjSBxTwPEruUHz6up4tR70E6eEO8ImSXQotbtt
zWoMG+0XhvUUNyRHGXnREaQc/wXzqGme9LFTx/52xx0t8BDYrsaI0CxFqtkHtDN8gS1T1iLSyJw4
nQKAbiHlowv5J/yHmaKzySHmw2O5apkReOeuzOrSxoaaR+D8d758HvLg0WaJc9zUe2cV7qeRkADV
WLuHLwJrFqCck7Lp91oAGVlGQXZpoK72iKfpahHz8GgXUU/tG4xkGbL5Tphhx/+AXU8PKIB3TQlh
H8SQReL9W1UXJEzA+Hp+wE/dzIOy2f1yZnzULZFfIlMA4m2s1c49VPpOvedidDPO/fIPR/1UBEwr
WPUe606/Xm9LZxjR539T/440z57MMQk/snx86S4Ztub2nL0XiBr2sbf+YW3dag04AdCe/SeF37G3
mNvi18RyTL/RwFweINOu/rxRFzNdZbyXiR23oIDXj78SnnmTXadTy6+SIRekEdV+xUAlVgxjqfGg
075QpWwu8Kndyj0qhZ/JKpEePuE65p0KbHPRKbRQcb/3dY8mIK8xUX0kG0PsYpERvKXf5mhY4wbN
Mwz2wvVvBRLaPHPV4f6sUHfNCoRnfSzTnCRzqsOkH7PTXFYVBD2/1SJw4B9ja4kJHs/3iLnDLuvC
b/H1JRJ5/ovRfrqFlx/IYS5deBaNk4FO/L4mUN1olawIapJ7mfYpDcn5pqhL9vZQOh6W4XwqNu3c
TfYd2E8rOq6qGrd5giC3hG3kBs9LZh4VJxSbdL+69a0XNlSEin7MpNsKkRERDvDDxGqyxykZfuBJ
vO3WLW5He+zr+Ui7NBZjL0DuM57yNXoebA39gZNqR1oBnCdlaB8shbL47Yx5zct1V3wE6M/DrOyE
m4ImLNC0srkVHj824ONhRJDCnCt4cDGnqWomALR5WQ2+rOu6WQIzRvS143L5d+yiO3gY0Eak0K3n
LMNCV8pjVE1wm3xjDNRNukcxCrJrOBBvk/ZMKdUAXq3VCwLe/1nHbrYF6X+DpQxxUdopHI4yfBC3
FnI2F148WosxzR0P+IQvePiYb7U/VT9Kk4jnGxLmMjcIDwI5pC4Y2GcQTNjFzZlsgdjejd2kw3lf
SAiSxBztrpp7qitDyUF9SwzYkmgJMxrZQk3QmBYaUtzw62uP7EheoOwrPaeKcSJFzE8NL9RKGK80
Mo7jXKAgxLl2UqFQsoLG6ZTOkx/lRl8Lt7VpM18fpAlqP1kC/KY2O7fl35E2g82VAY1fHVBEsKoV
lmrohSXcEaRUfgflcaWjNL7Vy/+Fnk+d3725HhLkDFhKElRbcNh7hyZWqxHx0m/beu2KUzxFwZTf
wImBuw7na9Ev7mi/N1PLkD3RvCs5MyjTrA3UD6Pl2uKkXRPxRwYAtRBP3kuJeZOe/1tv5a1es5My
58kWfkD04GKYldeBi0MevGBmEwuf9okfPlIFt+dlZ+D3VWhQy2DKIn793GOy9CepOJ2EBnddT9p5
lJJlxAXQB43NT8xK81hfJvL4zatSnppJKhnOIXxWMewpwqi72YMttMOpF4Rrw45TsveSb+UjK8QG
MnvZBOhUgZ0MPQrD92zSMEPEGd0InDXc8d30dxKtlFUfJKQXv7w4rA6p7rGEIBSq1j3e3lom8awH
cU4Sytm7Kl7wDGo85avRVTXIJ94wKnyaDGN/5zwZ9hOqTwg0iLtCKP2BTNbBk0Cm3Q2W/DpO0DAn
KIz0dc0zatsC0Qk96nMC0l7xF8CGVG0m8gsd1GMvoxmGrn7dsdxIeTlYEd3j4h8vXvPJQ/0kmbi1
jyWQw9WHTiNcTF/WrhMXeJqe2Gt9EHEjT3KtBmfUBR2/j5jdwRQ9itvi4hW0+MWQfIL3hkUsEI4s
ZXAflAfwH2Vp2f85h6Sc0bjztycxgyQBfN6BEHI6yES+AYn117L8hED8Zqm86pErkyYa1kkIDffP
kVdLh56blzglvvGx4MSXyKJl+hLOzIcWSPr/1qqjdGjTeF6XVNhmpEplWUDEOC6dw63ZwgwNWb/+
P1mHjpv5XBsSIcarAiVyTWovOjwTMX/M3hTA6oVr3ZJUbD4Qf2E48E2eEbiWDoekjAexyq0h+EGA
FEFCDCpo+a6WfBHdfPgvI6Tbzy43lxsxGIq2FsFhGgqsFpBnan5InKqI7/ubshwbwrTGqM8ikqLA
gRtJ3LsKDTj2q7dQGfHQK6xE9B+TakmhhvqyZTeWmxGfHent7aDTiBFi3BymJZhnFICBiQy1sWQ1
4YtviSj0OPUd+teJzBD9OPaPPZ95TyZcw7uS3Sftq7RlrWIybbW2vkWGDcVbeUtDkwoPk9Xpkyrf
UAhDLOl6ydmPXhK87MjGJdOzYrYhdMLv0Etblc4im8rex+80+YQ0XeDX+sehEDarxuRq71YwHmsd
PXzsD5mNJT/O9gFaJFL9afCTE9GGRErt6U+XIzW/lhaijzebNy6Yx1T/6VvkR47iYDl+JRhAEkhU
YLBKj8DLajpJg5qab+LrjXUK4gCU6js9Is2FGZvUgOIV+EHIw8L4m+KyrSZEP6UpcVHoqcEKirH9
O+KU9532pqU+VIvXfd3MnXHCks3NNIP3hpaV38Lmo/lhQZ9xghjVhHxm3SK4EurJLmqLHqx9ZCKE
qWuTy6wcZhKXRE1xdFOVqYl66Iqc+uw2UsOjeRrMepPrpnKYlWZyX/aq+wJDJwSzS/zhAIND4wGa
Wv0v1G0CUPkkuBTvCy9kFVZb553iC9B9IzBPCZSRvqHbZEf4dFGRtHkrzbzLZq0M583JYgRjn497
D2YGtfE+/cBiytXYA5LjDtU8ACIHcag8PjwpozSP4X15jjXBug85w2N/WMe5QT79y7EpX0MzyqjL
H9yDBloVa7kYhVP628i1d7Nt38OzMhbpSmUEAKGnEGB4B9QR6Zs0iQyR/yAognoljUBQjlGmMAMM
txcHKmrQ/fixIg2XutsdUbgp/JiqvXuDd3wM2/WaFKOvGD+3aMiheZRGHSdiuQpYQJxoaiEzQdt0
c6rdH/sVqZg5hKzbFCOjGJYlfTtNak3VYN4J3mF9zdjWLkmPA6CYCg3YEiu7hFF2NSBk1Pn1AR2V
x1NvDKYtYPFUD5SwlyilwJtjy94/fv5w6pfd0NJjlrbH8Up3DHoTDVL+ntfOdTIB8yyAawLsUPBK
fRSw14C6a4KBxLkWqmNmhcnJESKVbLqFqh84kPYD4DP9Q7roYiKctJ7OwAeZ/BsALhGF3SCpiwds
F6PKW3oH61Jq7njEAFFDbra7nce3Qs7OuDa6zz1Nciiv6N0sN4E2w+Vw2z8iN0BkAtqcFJDZDqpQ
XPb9/58gKXSFpS2kRfK65uWI0gWceq6AfKxiTM0sgf5JJBo41L83z4Y3P5Z64Zdoa1KjiRSlUApg
GHQ8zX25sypNt22xutYD/6szcsQTyyk0Ufj6+gR9rpXuJpKZpYt/eeCXUAQ6AnXhAIboo2/seftr
ijDhsiYvWdSNZ26N98FOaLsLCDPP9v/I4soiyAsJrQvJ28K8kCpHGLke6VwTohTXh2RbwkM7STLC
IVKSwyfZJk2fHQGr1FtPfCGCUlC8H3o1BwrPdwSSUqRBherJO2ytzEJp3Pxhog/TW5lu/dfvv4i8
HfyfK9bm7m06S0ZYII4/nExUfFWn/SfS0onSnCHHKaDl0qjzWQCZBhv02OYFXUV/+zhtOmIvSsfj
jwMDGmR8k9ElehSt4C5muLFnusdfdN9IRrU3+onRsruDWPv7X7MZ7xZS9fNGkSCBIDvfByDHo9Y6
7UEsftDQ3ak4yeom8GaikMBvubhj3AmZqE2tt1H6Aelgma8UonfmCeJ7Jm7VcD+auOjPhEdOtxQb
Uk12f2peGNtaD0SXqgahu2lFSLekd3+x9U47ddPDtrMuBcxsOWaywnFliyTP/4AJyP1/Wy3OtE90
VwYTzdBcoxu2kchjm/GRa8uuT6y2TaPoFWyJ+CpGv9qMuLMkQajIrJof3UjqX/wBgTo7cz8p/9Yh
P64C4wjYj6hIHN6hznIcPomxpyTNHhw0Yycs5nzXAlwPilyPp2wspF5fwgt2ilChxEeBybd1ROhH
GZKhFR9ry+egl7N4BqCVqggjn8hN3aVJjtkGDiItgMBgrlWzhmBOuU9vPP3yG40Bssi0iSKXY38y
S7KVjEOfD5nkdp0EdHucdszFIZDFDGuFJ7dUpE1l/9iaKMco0cVWkzV7+Imms3+24FunYVj2jhro
ErPsPpwh5f/zozUJ1E+apxENPS+qWU4LCbG4ZLdeOt8y8hRSmrLcVV/lrjwIKHFSIrj21ZVPPCtF
bofF+1ECtD6RzL0VxA82w9pd6rrZn4vi4zDrTOavRcZz67BV3+cKy6VmcD+vBka4sHgKHibtr3LS
f8IOFDWVGq97oZNe0N1fd7CB250s72EWU1W/8J9VP8Q4vUXZZzyktLaihHASmKXFfeMGn3F9cG6p
JAdY5lj9pXzlKpGrp8laMl0pWtBhYhvJYxIGJQI+KczAzQHOakJ0i8mqok99WK7mmDUKaswmwMvm
tTLeTFjM7+mGaNiXNcaeUp72uXq2RxBOgRuAZVvPxSX4QLwRB3FjrFwGfAERDYCYy5caFraQ/+h0
7J/qndoxxdHzGi8tPXuckyPQoNALYIWrZx1nYJJ9A9GjF2JiSy6fhlf9Drdlx6d7y79e0WTfdr6J
F1Jqo4Cl2nVzpIubGIO5eCxckTQTmizDyv7s62KKMtnE7w8Zd/VOfu9Lt2LtaWPIMvLqjbqne4td
OPPle8fNUaOB8nCJZzyzNP5iDjbPrDuIbNMCMeIxRKQkU+BqhivN8MTuCenOycjuLH88DP4elYKN
yKdns8FjkJSZucMJVWjUk+qWolHrLIT11LIjS9BRcPoywOQjS8HeSrJylaeUA09DL/L6BkCfJCS+
t4AIN5wFd6D8AO4eW2pV/KlUpXWc0juSYnu7tgU937Bw4c2hzQaRX+0R8HOQEjXuHHVrOOFk5Uqq
Tj5XXz/aZBDZ6beZGs0fJ1d2zWj/CzX3GHk+9MTCWrvFfn2GAykj6XKkRC62pDHp1TWuvpx0mowg
lnEP8KfrRGPtxcerBmt1rKsdfG4SiBl4r/A/5SQHGxdZdZPktbrju8SZ1zhem5gownBbQQGo0Dvc
VDydoONEMwT2DsJS7c4Jyx+Ib0qv3RqkDN8y1q0IUB6y9CvtrtZPNcxeZiAnyxGgpkNNWj31F3XT
C0whFbac6jmKsoQZknpMYYqUdvjFPNfmHsY8F3WeiJ9HMBoEs8rR0Y9HTu54Tw/Tk9qRYlYWbKV5
G2R8kdmvbIp8smrtZHJtBuaEdaW3yZELk0ziEhQ61RVrn9QeoBNEr7zyzZ6Fpg+B0GnOG/Ue+VYA
iKQdwfnQpOzbA8cuacJypGPwkLl8Sd93BOtUOCwut95CW6HuzN6H/D0o0D+LXFdLP/k+vEaY8DC0
sVtAXyDTjH6Z4lS1tgf6keukEA/kA6D22sX0S+ZoFMFWCYam3A5lVnUsloffEOdwjODzyXiTrIk1
9/yjSrjl7aSUcliM07mQ6BzPCMh5DqErTsixWCxSKOqw4za0sUgxiRlH1HiVUghHXPCuoaE4bLqB
9p2THaDx6cTBuS7gEfcS4Yx9l4PzDScf/gFzbL00bzmcU/wubXkzLRGbKSaExK9dfmlrf1pYNX6M
hY07xLiZq7Nw0SqzCcxTEq1EN8IKrbZhTTZrp+x5varuAFntHGl+ribfyzETZBi41jZAGbZw86/O
NElNvPb/XVaF1emmpcY9z7eVRrZcCtIF9kSvOPgh78FC1sC551GKm9hmnqN4XN4zaPoedLOVTBKP
U87Z3IHUqpWAjYd8n7CzkGWdWOblXaMBHH4y+AIo9ZH1UDQCCxeyGyn+tDBqOu4klvNUEv+KioiK
+RBPUt9GsrnyBSzSNV7SPeJDv9aaIpwdGbmMZ2jXGsGSZ39itTfMxd+5mglJ3Y79Z0h1X7p/2f3n
YvHOLY27x0aFpvtyJa202rLjcGE0wpOZJ0FGfcoxljZSkOTxAmOf6e635wRDhagy0Pd6FXS449Fn
JWfzMn+IJEOaeNz/EY1BVL/1+ZNRGHjkE+8y+SHydPor/kSCoYXJt4/2MriKjPrMw8VgCS8AHPsY
O5k7qYCBxVkRh3xCI6GjfHFszfuDPxDQAe/ozpGCGBviP3v7NhukFUD3xAUIjibLmwk0Rza2uAFY
faAUp4WnDJXcYhdqLLp9yFo2o/dgy05BSegENEua+o0kTtF2DX1EK7G3NJrT8WalDgcKaXBUX2VE
GpBtgqKiswaDiPLAr3aSZuCMeN+u970p9A5kqs6sQf5+2bkwUPraLD4f0ur6H2MyLyaCfBsyfbyX
mTDXp0MEqcxZ3G4lOG+ohaD0/5EX5Fh0/L26C0NlrLcQbEpfTUrJXv4IJMybEPth0Sg3v+Ha8e6c
nUmA5H5uk6KDht2bjxwEucOFKpBuxD1GDvX5o383WeqeKuEXFCipB12ONiJURlsb3uvjmorptJi2
muat0X2sDbAc7Ssrcje+Bpv/24GXm4UMf6NY1G0pw+yJ8Md4RN+X6yN4T1pyKANE9mxE9e/y5P34
CX5SSK0AiSldEtiudAuPuAvtPnZ8JFTcz/VMByjAUPn12nd1ds2rZ5auhgPSKVDSqQb4IoqjxocX
75aQNYVqPYvW5UuXY8m4QvWPpnjZGzwAs/5DMPA0gtr52/5ONmTCsiR7B//34KrM5IHV6YM/6K5f
WiwVvXxKFfKXucuPvniGBe2WkHV4iZCxPoArmQ57PDokrTbfQdBW0FJZUzTyWGXOVt59lGi0eFK2
xahAOc6blIIuz1RgNJu9breGZlu8qh3KpsIYDSkj+PgCbevjr4NVXUIsic6+L1rNItxMzuSQLjKM
z+YRrY1/VtwETxDbioXpWiniHE2nzErBy/o3Jdfv3PsKv7otW04tvk2LhorYZ2H6yAYS+eJwFtct
C27zPFbV0cuQIfHznXYvexwS/o+f/pB+JG0kEIiM3KuOvrfQH6SzCl+pB6I/aLyjCOfFdUOo2mkq
GkBsHP4uLLPBhtvd7wfz3ipth7Clg0fxvG+QFB7Ho1WtIL/qegbCto5pGx2c1NGjk1HFlIbhPG40
Ec6rsD3Oy2Q0FxV8ItzkOniCL4GfOc8U7r3F1OHhnAtyardL5MmxYScA5Ml+7dkSfW8j1uUhgUGP
yX5r0MAPkszjcPqylFkb/zWNxzDYxLA3leoGRqWGriAKaCx6ACwxYjcArw0MuujlXP1686u2lMn8
92eDH+zw91o8Wa47i39N8cafkpZWI34b4icxCyT+M1QGJGs+41lX0XLqruDULOHogfJA8Qt/2AcB
Ffm2pCPy/UDko89l5PDTAWx07pxmtxExN9uuJ2TlIyiQfRwmYWp96Nvy+LvMSMA0Oeyz+O3GgPKz
5eD44x6qbqXU4MUW0a1CE84CoyxaCkBoXf/VvhxXrz9bLup9+nnbBnxxXd24uXstqacB3cU+yh/L
M7jAzA/bzbFgrjy9dUBGGLfApKT8b1okgPK8ZiMeAKVCfTfqAlF4d/LwlyIpFGRmoJLasyHG6X5E
tRil8zJU+dZeWz6RC8w2Jc6a9IGJBa2vnO0guRGRWZ5gUHGAqALy3e3eKReKMiarsbRx1xnhqysk
1hjQYBBG6x06Bv2ksj1p2RM7UBCcBEPvpzsjJhk1XZcURpt6MyH+dVwqToIJQ54UzOBsro4JoBSo
+N28+vOHltaWz+OGRds5RWPIo5n/938MM/tBWyqZd+IAPIAZpjWjI+1pGqqTV5BGApFseCHQ3l47
m5kzeNtfJTM0XrXcceLNhDApRP7TTyrSH9irtdMxNFqsjkouEQR9bQF3WKIjQZGxNayhv53Ma0XM
ti8tTf10yU4fPMgi3JNKYeWKBvdCUdgkvXikl2ps9ioADxgFNbF7KrazWUuVCSMt5hcO2cCtB5yQ
m6MeDqyHvB2Egt8+IOUOJP1+EZcYdgCm7omfLafExy1L1m5fsewohWBRPkt93yIr2epuap8tOVym
NxBzNYOJBGIqxkcKUXXQOepwKgFI86934tHGo6JF84np4eSFDlzbOi6IwUDoqtJGVKhvn2TpH/iv
S7p8n5kEapIUhKhIRKdwOQRtrKoDpH71NK3Jo8qcG4YUMYW2LB4L5v/PML4LYk0T6A6oNeniVWO/
DZAmmDH//l7fyxCCk5bGzn1T/p4UEei8Fb3oqwcmQS7c7ARBeJdlhFj2eWkwJHf82mvX9eYi0b7P
Msyx+LIecoWiBEwjGmwTCmM8B+WqYEXgBqijQa3wD+7V95YtPw3IMWoT6R2Fw2TZhiOCQRrumWoK
3sevlrSPwfiU2yVnRTU9vIAEOIJHR33z2PFgjU2tLp/8O6MXstQ+Avo4AV7aSlRmIqiVMbPSQprw
M61vPq7Mt1uIzGIRgGk69Td7fS7WTZxspajdbyU1kVXCahUBt+flT1BPEO5TFdyxB0/4FXltdBtu
vpo7q7Rz1APwemLuNHi4ybS3+oeCB/WGOXlZv9NdtuhY4BFjG3vwtYApAgKH0DIHrvw55EVPJ67M
JnQBmFHTFiZYIGki6OboWj6VaMiLIrebNaH8NFBldFw09tJvrvK/FKlZ4nS6KK/2HmUn46ZfbHlo
kxwc8vYQFo2XXLVXPGSWhAzU4P+TauopRHqCu+A+BmOR/aHEhhfQ5xBT2MeA6HU+ub6gJtL8WYw2
K+iNx1cUaqR8OnDpzY4ZIuP/O7r6GnStglX4vNr3g07J0BW5gsXRPrA0XjVNJa7yJTf+LJm6qozd
CER/ePNXQ/lJQbVGWec+TqWGiaPzlF9z6rjUF0+EhlKBOrZjVNYpLsn2BrPHfcwo5AL3U3xT413Y
/7kf0jFbw5l0K0jyPklMEWdq7fYuBmNcYNMHv5NNIHiX6RTgTc/5oDr4bSPyHWpw7YvBGdqxBYxp
wimDnr4XeYxTAwCrUtQ0RZhnIHjKULbQOodNvBtuOoW8b7egFwuWs5qElJOu20cmaXpN08dXHzpw
YsqZYdviTD7wunv9ZRFrk7PIVuC69gxQ4IVW8WOteGp0XiKEmeniFEpc0f1O8g8D1MrJyRk1yJYA
jj57XrFFHom0zQR8UXQ2BTZmrTRvj8FKrA1oL4nkAyUgJFzvjuPnjrdbLDZIrbWGxtKo+USncuPq
vPwIsjY9XoL0VU6BYA+X5Pxpyz1e41qKAPJP2CO/vrCTwQMK96BaR4XWlSejw7rc6jKpDMRRk/J7
ga7PuAGnBcG/7ufrfdubHLFTkj1dqeSfwSmQHpNmQJPGovcrp8hoi4zCzwkKcQQav20YTMiwAHIy
aSJRmmqtAQzQeEx8DajSlxPpnikil0Hxk6I0gzGlRHfzZd700HiEYZAX8k+o8r8zqhevSw8ogTiF
yJstsSZyNqVExCELREIS+OSvyOg1TQjR/Ag9LHVtfd0bv0ZlZR3NcozMWPCQYL79ImFufPxa/1kz
VI3b9LBrzH17xPCCYJDrq/XlOaMElr3VtSjL2BM8Aqxzmvw5Lq6YitgiGQfozfwjJj+vczBX507t
kwxUlNqetlsW39EGwDDRBUWgW9eMsFWaEUKQ9OWuEYu77nZcHgRgvbuIlZW0nGgTidBh+50ggkuF
A+N2YxPmJy7MuvvIzFvKaolPYqf1N6CTQ6a5PQuLXfpCCdUsf2PvfK1fw3vFFL+qZjK4vtORIc8v
oCe/EyPvV5c4a1Z7O1Jl13gpTSIFVjsC75k4kZ1m5g0iiQC6ejU7kN/SUYnpgVfSX9FAwlB35M4Q
5tlmV9TeoVsseD5eBnT/kM5aBNuFHoRKCrPzcYjZAVvC2x81CHCPrPxAAql2s9lYZx3VirYwP9s4
o/VNV8sbBlqkkL0cp+SN5+d7A/j3DMTsKn/aQawOjunQ2VKQY1NtInMWavD8qRJQg7z64p5HI8sL
fYpRVGVeJxDF0YRJe84YkkMD3nVNrC2Csl5YWhJybB02rMGfqp6p/Ui5rlmuWbkRWAEEkNhAYsuw
+xQWRsNE9xxiJ0T1EWpn64ESIJ+5zv3S0WngFAAe+YvFDe4icYmrjFzaTh079ymKgp8FLNqbutaZ
L17vfYhTpryR43Qn1LTXgR4K8gnrpBNdAZ4EC8b92pNBz0tLptODr714SVEQZURfVz9YHBpUbpL3
H+g9FNL8PEAFerTMpfLKzPH8qBp7Q8Why55nMIdmHYlCgWGSbsxrCzoTMG5vikbrsyqnb9Pn0MEY
3gGuWanOsJjrQPLOnrnroWP3QHYxrUDmAt7v8NaVyf85KfDQg4yHkpZXUgT76olug3aoKQsYauqK
9lu/wgREFleGlXNgtQ9mJJbkQbuIPYNgn6zHyMjpy8qm9AEZVYcaKu63hCxQp7ZYOVqZLb9oIj73
tPH68LspLT9rtwTQZOPFtwPQSRdA8mPHvtiriCLQC8e/m2wdcXpqu57r04w9wqdlNfN+DcwD0xeM
xbanJs4ehrNvqUDhIXCjmZLIOy8gK0EIuU70t+v69HGvGofTFM4k4NZfwuaHiHUUqNsIMOmSBgr2
LONWbjs1ptEHOiJRu7Ud/b2TizV21bKtR/ALBhPNE1zELKoAzK+h/SVYNWdQfNztsQfnpYOdavw8
Tv0zwJ2AvVNwYqlW6r34zg2JIAGxPB3E4p8MJP0A6RwsvgaYLuQaelZvTStrQEr1kRwc4gHf2+P6
VBqt6bpU8GpW52dKv4rdS4j5/WOm5HxoQmywJ5TWthITR01S0FpTi5aYNECfcaRrUCSTwb0gY4xj
vJ6xSZ2uFnYx4e6nFU+i0Gr/jGZ+cDxSoqVArteF581Zm39pYLX9ZhLCDI+K9g9jdeJWKsFyE9Xb
BBsjxAr2r71F6A9Q98Y79N8zZtkP9gLEydioKExYwWthqwcQ3tj0tXiylmzMPM8AU+fM2mg/zW/6
u8VZpKRbqnxQHq5kfnh/UAcevWxFXmEZqabFg3z4ej5DPxwE/UIsKgq7OdzFi7t8DafiGdu4xyeX
UXNcLEQBCY6tkJngNtmTa7bL5TnSFtw5KiYT9FvudDS+aRb8D+aVTQPfeySgUet+CorHvrUPw4uN
b4gOsOr/hctV5MAG6zTM5mzetCbQPJkqQUiZkXl2SUd6XB1cNEAaLQup02+BnLPUNqjtYPV2nAbU
wIrdUxftfo6kTpcTYx8Zy0ab6hIhXOz9x1daf5tbQFvRHx91OF3ct54ObV/zufUPOurrheSrIhPE
md+7jp6nergoK5hr8wSvh8wI0UTC0v3GZpA4YHOm4WKwDR5xn89QKwzf5Ycx3HjcgEXiui7VKBOP
PNe3ePAOkvDDjFrU08a3P9qQhsgT3wjIGROY4GJ7PAzeaeASXhjnrgIuZrfUWEO+Y6kRhzN8z//1
5A6VbeThvRXLdmGTf4ZdPhmCuygixrahVqO1UfAwQjKxFv0q8PXgLDyVSceApt2163uWIgpp/eWl
FpSM+i0KhUrEhGm9iuf2xb2y1gxas0cUQDc2JAeGgLjXO03rg+89CxDcDsrndqselSy3hPWqIg9g
YZdtsXhjun/KcuDT+3ohfR1fIUabo4d2/YqRF8NscoK157TT/KR15reNz4OhxLGXj7VNx5Wbx12V
mksIav33+iClZtpGScwsitSya8NZfy8ul9Z7DlqfD4b+w2ANvSep398f7q4m3UflU+rx4RvcCTD8
GfN3HGv58GkVm9xEHoY5LGgTOGgFAINywY/pnpPu2pL4sBjumzT0Ykh6nHxgIHZgcWdOXlRwSU+f
z9uAJzCQpluMHw3ZmiELqbWGFvAhzY7N2DKsSDYgYS7uz/gIicc6F58uzBoLhs3Wd5lpVuNZ9Hvk
W4Syv0ITx8dvVe9Mar8Pi38O5uu8vh3vLCSPrOAUJ2qmLvokbZqeBmrS+bElU/7PP60F54C5kaVT
7p2HhJgWiboKBRBZOYWnvIBg/MbBVNBdLSwX4JI/e/LbsMEHQc511Ryxa7ZwMLIcY2CD+YsCVeoR
HYLu0NqjPJnB1NT4wXhKE6O1RORRaWIwGpIj9FSvTz+LFDURwCEBOHsUDgGW1L19kEMl0GK7MlwB
yzAba9ajhoNYoNjVhm4HxWS2n9P12WbepfLch366hPbdaQ06if1wLrAHWCXik9Zs0RlBCEbQ7LFy
mOvRfutsHf9wRC5MQ7i2R0u7CvMeHOMJNblqx0EpNhgiQLWCQtygpQn523fITIO2TJFhWb61EGGj
3kUZojLaJCSB14tGhK7cv2Z6ms5R72g3HFhdeqVhUUr10FeJ0zs/Go6+PC8HtcUYz5hQAu67w3FN
sWonYOv+6nn2tpTPEnglonP5AIHF0ca0BRi4tb6MfzmxCLHPpJu5KgRUb5hknXeh9dKMuhX9+hse
dW3hYFl4T1CLHOXPEms6A4H7Gu8XHqkOypM9uZK2iMelYA947hXptm7WezFddLaAYTOIhyI4biQZ
u0aXLb7pLGbvsAtU4Bm1OdWXz4fNCjbwBK4TN5xgBcpi42Iff+C+YHZNqXCMPN8ZcYsfGnWFiNZx
S/3wTC7a5KhJxpefNEol1eB5GejouLgqwfNz4Uq7EIphCvIRrrAAQRvKj7paM8gv7/5TxkFkceqW
lOPqzod0Yg7/vyOuju/wD2ffnWcCU7+3jx+eIpNO7SBUQXRa5yU7EJuhEr3nQ+IAg0dvACPbz0OH
6LZsP0G/nuQFBp6AxPLmsu4rt58B6DM+RILgjHznm5fjlIuD1WpB7X2ekr6VMUY17fBAnY1g/416
ohPGkGlTYCxycZu1qAVg3nF4wf7PJ2V2T740SKuZfsfrqWtvQCZISvUduJAG7zb3fubtBwio2MQQ
SMmhIld0zwbTwIihvv6ybBZUyr+p9pf8OLCQMvsHoQZzb/eWLLilLX7P12EBMhDh32KvP+dEmqoF
67J5NdV8ERPXMEabxe2mU8uJpUzrdZBbdzBSLKbG48RT7su4eAE9MM6O5q5EU1e7rvhe+8eJ7gbX
JUddYBt+OmfviFVVST3Rm4mklkEHnS6dlP57ucK8CxTTzyqLqkFcBORZV/Na2U3HUSngrwCNyxu/
vCLW2+WtzQRsKL55/avEFn6MiDPDKbWV8hesnXIDOg+0cmtox+nnRycf5yq2vrj9zdy2bylfPeAO
u0phL677EbjhsmlXzUEPBXz+q1N6TRsvQwTHQZ9nAY+gmLSGvsdV1Ih+YkhDXzuoRhbTo+MA/wni
PeAtFIaMN65zU0cCuSKCk0yYeUxc9sotRFbN8WmTZgs2oOb6KjIm7cQHXFXK2KfnkW0ScPHO31mW
qqgv4Xh8CYVkeXNqg7/DQ3T2386F3e2zM64utNbNkFKdjc7E5r+1qEyscNxXFtpo2+EwB6V66t5Z
FBzadK5wfitcGJq9Ydv4YS6+WUh7ugQTAGXwGhVLiE3UBMfwY+HmeIuIIY6npbl5TklIZBbRSJf7
NU2BQJqmVaD/EiMDDFbXITx5TS31BdzWyTORylX5m+kPYS0SNSWKmv3CYfdrL8jP+xp/weIoWTBV
8Csd5xO8Vrky1Ioc+hnK2Xr0TrVsaiZLddnd6pE7igljxBWkNmJuffOo+e2LMtp+4pTXbO6KeXXc
UprVFmU2lEqeXnewhLaUjCUGZrF7lce0vebarCKtj8dnvSIStmCcu5iWbLHTeY0yCAcZ94cO8o18
SeA3+ymfwyylhYhkixlyeNBwyVmOQfluqJN3gk+pRHhfmLJ7iD+q2vrJzTNH9eudrJUyE5N03Dij
Pv1OFEhKBN3HCzDEUzOEffcKCVcIij+51N+VctQLEnGCpOsIabYIh5xnrXuiR9ZXuVxazKla4l1U
IPvvoiuEo+vspn7COEAm7Iq9M4JM2Dv5YrcQ49vyaWDvZWPSZPM1d3oOUjFTQutZwEs4uUVNU5nj
UUcv7Le3qk/WhzDzHUxg0MyXYh8JI58YKGGCno+xAxLhxRqjjnAI/vSvjNDZkwlev7h96pkJy2DO
I3jozdAAe7E/W5gcKOAurFYHulsZx17UTcQ2ATtTo4FxL9oV3jlRaYHYxkAJhB7VIiKoVSuCLsNV
Bn7HGAxrW0ac6fuT+JWNGK6nZjGD+jPaog0945Gc/eDH5Y8lhsVvP6jGt5FqrjnNjwCbP7R/g6B5
jgnAEYi4VN1hhEMjidGkP2BVz2f/EPIxPaYucUEbaeVvzWMoc1JJ+fypUse5Ml7NMFYKVnKnuzhv
OXb+RZOhUiEmyk6lSA1QBRs3/sWdrgfka3VwMkNfvoNBvQY2ra/ZGXlq54rmk9CZrd23ASXM+A53
19poDFvUE4/PDpn/EJ06bmwB6AI0At1e7yPTCM9L09XT/myhKPduFM8vHlIyCY182wkg0AQb5g0S
jvK+F2DhzjFb1AeLN81HYRWznH4VAplL6tXp5b+cnl3fzWuaGzOv8ePBhZmt/MIYHdKYjsNOJ5FB
rPs1OTq7ww9Il2wR8ESW77woylfX8bDUCsClFMfu5U2mqsAC5vRIlNQ+bEPdN8omxo4knDTtdh43
w948hxlDNL33SalKMTKjO/lXVN9R3PQyu58pGkJ/bdmOxKoHtxBPwLP8s1YjR+FAXc35M350lzys
6bHHhS2GL19PhBPDop8MZc6HD6zgPAXbBwjE5rzj//z0o/ovZHv3Gc658OMEgUwq1I6C04yU+GUX
Yo2T4wiPEVjxjTVV3BqgeO+6TayEAE6m5oBqr48hEV5urh3hDwM17hkxdN0kza07vaXqOcNmGdTM
DXh5B2lUM/Fx5YOUyX1/VbWEciHR6ChPvr4REOHIJB5/Z9B40dIBrlASig+r1QsqrdbqOtApwp8a
YCqNjR6x3cvEncf8TlfinwC4K8KNo3+2/G7v0dVeJTevkYKriGTaw/O0RvJM6KpIXRvam6XZ2nke
WKAZo5uuI9+21UXweELZbsoqbcJLmrtHvF/CgnyllkCrqHj6N38GOlEk1FvBtB0q6oF9Xg8snpOS
Du+TY7kvD97Qsfl5zsb2BGSZB8Q/MMRtrT82cpVoGzpY7GoKdT45o2Je1hIr1sHyWPgTSbKCm+Mk
NeX/tKrKZAwdeNY0K1QAVv9wi47cUi5KgNGEGakWYIl6c1sx6hUaLh8F18GjK+9JqBOKkO5rNKq6
1UyldNRimIb0BtIG8K/rOWC6mQzsVDTvbziyW4IwYPt/x4FuPXiLmnzFtR+OsLrA4WniXr2zOk6G
AXPyuw23H2UUyyyqWsbxT+XR0KzAmw2Q+4GNnLeHtb+QxzSSUtnFDm+gFNebyOkw+UdxNd4p2Y9C
ywR4R1I2ZPA2gdmIkhfMLgEtoOS2YRMukrpzvdReHphzr3JXo0eM7Jm1znDle3s05vLoLZJufCNh
Rzpo3E6slZ8fO25aAAWy8bCIWiWKjd0gcSAJbD1UjlGIQp1ItREZ/YqQ6gKVuNFWsyfaNsmrZ2ym
Qkemw+5RX/T/fNWbk42Fbhxlg3NZSqrF2/b2WVsuoF1nBxWEqyGFK/bq+pjw6YUhzNcFOx9SGwht
RR65lMnggPaG7MZ4iXPRGDDcwNx71vI+7JPhhCbhHbrlT4U2jaUWbIEGNljWaMEXjChRSRxG+tHO
Hlyi49HvJm4uFoQWzNMs/Qw3t7eezjaUWn280bnNGITjhBNWYk5u90pJQ3vi5IjQVV6BPO653zHI
hwo+cKWz2Ft81A1jbd73ay+TBsvPJmJNGq8vvoAeSOzSsE7fS42LK6ULe8H7414D81T3CRUnOKLo
/qwsqyLVEQvWS7drDNV/Oow/9LZFpVf+3pXMScgs3VX6I7DCOAQYRjEpSt5NrnQTfNs4P/ZRWOcf
o1Of8grvojlK8H+hvlXTocEbsCVwN1Qd0DIb1qD8+7zmxgBqdq7U6+ihBm68k+QUMuADD1t48KHs
4YhPClRhFal0TSOJUId3yym3hVwZUwLDE3H1NieKHytvBh14YLzFf2+FZxwH0ps76KDP6tzye20o
qC4isR8LSPTsltjR3nGQiY7VK1dOc3klrn1xwybao57Kt3wzIwvpKvvPBp+lQTSQ8hVdZ+DvbIwq
KuM8gpm/6szkabNBIvvGFKUgQ3Iig7QR8rk+vgmlWBFQdPDwUUNsichkekLZ7jYCfD/BrCTx2qYD
drRl40B9nwvxer7eAy8CuAfv4rbFHCGVKi6ixccGVNOTp+9O8TFnPDTuwP6KIE+9eVllwUmI2lPs
KQenkB49t5wm7e6RwuKzHJbumNxH22qrJFP7EqxeE3sXfJcS1tOL0GcopTE3/dshUENy262SDtWQ
Mykvv5o8oWdbXS86ygxMEiZMXSYYgmB4pVbtyb33l6IkI50gE0TamrfpkUik5VfItiXwYsv+cCiW
X98HxrP0PbAQAGJsMuqzXJXAW/D3oCQQ7SKVZcJbY0WZchHGTeWFYazOisM3MjHWd6WcYjq/R7Co
G7RxZ7miAd+aYFNLRyeOGyYVURTbtG8ROTpEmB4CINdsWsIyMsmJgg2fzf+E8WwPo85BQhQlXV4I
ttLPNp09WQXRr9xy6lA6uxW6l5mK11ssOzLmg8zEX6+yWKYDfxru4a0zPdpQ1QdS6mC/6AugzpSF
ZVxQfDZ/UxmIoki3FFXMhYacEg/SPremZU/WgsspuaNSggdWmCHqIPzrKFe9PlXK8VYaBwSlLFN9
NQs56TUhrO7ShpYU4ERNPLrx1mbRjJdQiypD+iUbzGxmN5NsMIYGzrEEpMOgqnJNjH+EKAHASywz
QnZdoxb4RlU7FhXYxrtZWXFpIOlTK797GbBbnW9iWP1YmHsas+mMIjRwVjuDq/QTE0fyCGOUUA9j
EOhKGAeWE3/7r+Skk8580zhDDohl0zn63T8vL90sSHGmb5u5NdeCw7cWizTV9gTQaGvZZBKiMMai
+bs2QsZoC0f4e+BjvDrBSK+wRWxlvhBFVuWKEpqP8jXUQDompoG/wY7MjIpQ1eHJkFG1rB6iEZhU
cfFo3eDprLMqhDhkPR3Y+ami236PLa5I8qqt07MOo3c9rUQ0AYRVn9jednpaKfcWJ2iikU+fn6Pd
LfpANzlTpcehb8mcWumn86+1fNcTBH7IIx0QYBGrVd22s7McMcvP1LRWLgwACR6k08QsN9KLQ1h2
rsjnnurrMVBgi0cB78etysJhozXiGYL6aqQzNhADIo5SiHR2NSNJfmbNd4jPE7BUgwxw/QL3KR/5
BgEqG+zCzKbOnq5Gb7qITJbv1T8WBIgBgDW7cabkegBGjI/EviwPd61FOLf7gHbrKV2g8fdK8PfJ
XUOq1/sZaZ0AOX0flQwEZxMGyzQqCqvBD1daP7qLqmQWUaGMrvKKDgfsiJen1Qe6sLmzr1xhUt0A
xmGZ6EHxt3taDvsoOTb6RW84aJQoIpWnTnPVkhjswpha4xsPBemDJc3gA+6bsiRyae7S0sI0f51Z
h7tmbaUQrWErM7ihheXP3YdlrYlsy1B3ObDB/xfW1TvFQeMtAMT9vNzseyE3xMjVUwmqTymOpbRf
VqGNxpGZmU2JCFmPPkMOvU3LQxzu2tMOw1bM64CWeBFWYKv3sKphbWp51ZNSfWkb1stQYHmO7i1s
GRDEYpqfEG87OOyvTgcaa2yB24Um4TwBZM1agh/6eK+gVZPipkvQ8KBKaVfGwSR0EWYQG4eIeaV2
1TlaW9UTAmQgHo5cKW7FC92SIGB7aSQqZ45lN+vWxAgM+l+TiSReGO3rjep5z/aJDB9ee5cXJyK1
7viluus/QmwmXweq4f0my0fX8wsuH4mrzqPDQYRH1Lmtgwj39CQEv59/luvCy9v2YZu0KjVRq+N5
K8a5s+zWoKLd9vaB89x88vsbjPLAYEGczmbAx8r35du6GOKfZa4FzTlAttZHrbwO5sh7A2yeefbx
TGAHyI31Y4WLciZTiA1GXBpEHo4DJWleyjPOaSUeZWjLJoLDrE6u5BsPRGwk2LlJdDON15Ldn9d5
v9qSDG/hFCAlBBER5EhJZwOJsuxmhJSf9oSpog5imTCkJenkvSBkX29V2ZiSFKbdRnfWb7I3t/JR
QWgduwdP8E4S0rI3iqU5Kz3GMiRnXi5AoS3XbcK9AjKcH5zm5ImyWQcZEz3VSS6hb0B0w1joCqjc
dXAZghCbXyWu5qKVwO7JgbVy+DEIPe3/wTiUYJ8nfIswhJZB66xu2zOoYKfxJBDQyVkyId4wiacg
/pewyNe/0lIoZpZtqdyAjf/DL9JguyT2w3w0ny14DxbWl1lvtqPx5gXblfJbCv4KS5OWo0kCEMTT
yZrxZDnxQRnmhAlNbsBJabCrxeWCvxS/RktCnXBMbz3V2txwNlO8PcNt+OM81qPspPKnVKn+HWh+
cQ41EP1zVJkH0ThSHJc9bmn9tWOUibzYhaO6HJYqJPUOtt1zPtUxXEIDIKQUyUYbSS86hW1sKiak
7q4RGTh8JG4y+x18s3EJLwZVjGVtXUUW586XlGTKyRzVUBaXwpggNHAEHrgxhL7dRs02zz8/epRD
OsEBIKe8A/KBpwGwrIIrHAJD/dDTlmSqpgfvyfyGiYVbbsiJx08XAtR4fFeQ2tc9+j4fOev2ef6W
5GxKTLjV237I5ZKxrqgTCH0jTExGviCMSKWGJ60Ua9bWJjOkCtc24uTbtUK+bxSyjGqSqjzDkmnW
Xq80UbaoKWHJDqxg2TIqMSwt8Aw6vvrfUU1aaDUsC9X/2Te8WgclJzzry/U/1iiCHQ/vp3upNees
nPgGc0m/P76UrOE5VKPn+IAjm5D5Hvkvpid/wun28gfQgT3Vm1dkX/ZOunIveqgTY3799UFC7nXT
R9NAAlZOsGgNx2S718CjlJLrK1E/MrhalqyKl/KaRNjIpNa7I1do1qK8giH9OaoSNcMJ0/LzFoLP
CRdrifgPZ30kqB1kH7C8jbe2L8zjOPiY/+8zvNCtO6eR1hHdIDQl4P+bE0adGlGVn3Fv9I2pSGxL
tnQ+6TVOJjZFHdBZb+I48SzDSGwx1O9GNLzR4i8tc6R6hAq+9kOjGrXPyZYoSGY8E/yKJjflNPuA
j1F4A+Zdc9XA5k2RjYDRQyBJrlKqqgUPpw1FywGsBzJLVt5iyEaOpeT7qCNZNdRvei22azHtcvSL
8LR6Yyy4xJCmuZ9jho05EtvrZLlM27THwgWcdaYTlqKdawbiBE47mVMNGUP50dMKCfv1zbJfMatk
M5QDaPxKhjusyHBRQofjvXmWGr54gWGm+4SeK/afg6b6obn0MeUYn274RTB9z/94LID2cvvzLYUH
V7cz2guEegdeXfyM1IVLGNQypTpyWAfMLfstM4D3rrSv2QHhDQ89/2N8sztMHC5LZQ7C+vKOI1eo
hm5TdNlw2HDtIxy57J3xJLOExa5IKh4OT/TTZNcg9KDsF0k1+0pYHfFOdgv4G1msi9L7dtSvx+gA
1JVvIyyJ0JZo4X76WPaql3u89j23td/fK1BwylqbcCFTKLcGeB3KSXdbaMFVD1e0FOKEpXooCbPO
TDj3Y18I3WmAr3MlhlQDQhD2Y5xEQfJ6i8gUGOzN4n75Vv27y1DN9VM4Zwkk89UKzeJIPbUGho83
LXOyXYBJ8ZQJcskx0TVTSludscp12JpTTM3EB5E5ALl1tF6mVELAzhU1B3uZ/eJdyY6hy0SOH3pe
y2gNGQ+eSTtygCleMn4zy/sahkfFr5pgtxfGvW25fA52QzmRPYZzilKKI4K1CDOV/BQkv2JnkU7D
ihHEmSU6pqrsqgspN3deXvoYktHX17/pSXc8m1ZHZZF2Hct5XfW9vMeIMdpjUKXP4WeaHcIn+hSy
4vFML/SspYGQ35uKpG/fKVkTr4w07hsgUZMM4KDlQ+Tg19rZJRNioV98JEwx/yNwJQ7yy8rvmxte
aRtBeB4fsxcaigT/Ki/0QT5nxOjJXuuQfer5QNGFdQ61y9eHWWpv3ec4jAP5YEw5OPUJA21wtYrk
o8jgqC3twBNOoCi96pGz/PQjjQ1sLpwqVKmBTYkaBzt/SrK/e44ameFiohvhxdS99EyGZxYi6XKI
1n9+i921WEASc97ef6KJgKwpSeBS7iWHi3XBqcZosED7nyf0IVE3CAAZtmnAW5rjuh4KmnK4iRyJ
zzkcMSDuzEMkVHj5sNDlJvy1j0rbu2ZPVIi+Ty/oOVz1rR3VrB7Y3mxgV1dHz7JNOMbbiBdm+Tkz
CJAFJ++Ih8gyAq43B2fEX0APoWhefCYUYdSR9xoDSpuTykl9r8e8WVdPqSaABSgQXuQ7PMDEtrRz
lmycdNmg+wlGa6MUwKwUntzxIP302kScTppRH6z/wiUCWh+ALeYA/vudZmJhDn+ORiFjA9V2jBJ2
ZzqJnK1WQB97yRgsGLTbNIwhEm7sOFzO8rpdXps8Xw6OGJj6Oz4JlV7qZPchZxYD5fyGY1qBCDEB
jHipwZ3umiLIP7OeUu1efH24/W2WvYTwv/bz8llOfSSIHypocwK9I9g5g9VW3BiUTNYDpe/P5+ha
k/qXuljhWvlr5r1XRw3NFpvhGLnl+vTqbntbsUX+4OnwdPgg4KP2Te+Z/DgUJGWDPBHj720+NDXi
EVp1xYqNI+/PW72jNy8a58655lDWBQTtZiiRiCQBgCGWxSYdTXm8atv9otiQGShOijxb54ftKBg7
qcBAhceMl4Vc3P/9vhGzxgKTpjYRdPBSAHNzQCgN+GHLx7PsUGZcOepCfPT0bszTQspzXhGR+vkJ
XM6EEzgNWtBpenvf8qn/5kIemGu78ADJ8Ufvu2457royKR4fHBB+xc8RhO4++8wjmi2FCELVXPiB
MF50sL5CoSjnDGPzxedG1lou5UZB58bXtNyGrHLphBaNVo9SbnnIcTqaj6WIs29UoYsb/1tB9t7T
ES1bF+r/+cIQvQnG0u8HUPh2vLGMFhJnUhX95w1w2vDgrzpvH/MYYwdspQhuoRP2ifKE3yw2UVY6
XrhiQLHMKF81eOz3bv7X9pf09wpXYTRjMGacxy5zwn9a4Atc+RoO+oYrh4C1WfDXikeq+3yeAab0
RlVcWzPzzsT/HcIwhl19+4xKJVdW9eYL5nMUitQNhuFlyWsJ1b1KmtqCQqEZPScwmZjPYsRqU9Y2
poPV5ZVgn6oUQWIyvZj94vD1FYjY2AtAo+joTqXHXWmyTdyUkQf622Ixq0mUUwJzjc8EQrMJwBvs
0QzvtLUaTDgE11OI0XIbXzboP7jyzqnqcGIZyB/NcpyIcdcid5ZuWepDDoO3hsSDlJx1BW/hkySf
JzhS04ktMOVGM/KRrHyGb15WJ2eePOIchejglBBh9GiRSLX1IYW9bWjkFRwzN2cEg/P7AuqEQh3b
SpneBpwB22ZQa1dzgFtA3GklZulBuCazRC2oz8sC2b7sZSTlW4w3s6nzNBVkMxs/+9AuDXK2sAR8
j0GrHO8k4tBk1yn+bC+TdnbNk8ngC8QIP9DMikQ00jxodMVkrn8/2UMRe8BW8o49xTJULZwka8HW
cmYE8zCREkugnHVP1ur/srkGTtcFatrxx3iK7oOiI8OErO0YO1eb9SC7qpciFmfRNxn3eSengXuq
UmaWo4rIS81T18PsbqsoYD10nO5gMTLKFq4JAvVsubYa2tYVkloMbVRVlSWQg2TudG0Zq+HpckfI
oxy3/TmzNATYi5hW2mNICrtLBzaWetKwybJyPUHsDyDdjb1DPMyWMAPmIAQbPeCA2h2dzogOkna7
jyXmGkNXwx1ZLbFib/XaLxVbuYJdHB1WFHZwKxf8ycrpvNNSy0mQX+kKzD2V50PTrvw2CYDcXDFN
I8nPRzEcK00mSs0VPkc3GeBxRouDiEqVo5Vr6eEH30IIx0Qb9ua7U+TyhLX6jNESONGI+OfhwrFV
b4oLJfiS7tG+isEabdtuGDztFAfoMAaJEUZia8MYq3jCIRvICfbuG1/sc+Y9TiMMvrpfO78Suoud
VMDmRWRwtbw0eBzDSZKa/EVbqxBRwOS6JCHr+cLvLx7VWBXgZW+egpX8onmzZOXDmUgzGfLbPR/O
jCaAa+hD+erZNk/mbPV0nZ1gH08aBB9Jil2wVh4SX9fVlDY9r4E0Dw7wAOVO4whfpckcVHnIJ0Kw
Tymu44zge9/2uN0JW8AxT7K7+mDSNYBgh65v91wdN+aKezk2juHFPMC2lgXrfMsTYJfQNdsff58Y
6vmYCyUVAJQa3Yyb1iG8Ab8YzvXQ2AimPlLC6OWJsf3hDwM2Qfsva7mcjlXBvHuRSX9mEOY6RoHr
frIxD+z2iE63//dfPHlJrhPbty3C+UKtCIa/Ylwo8MmZ0709Q/LojL/rRw7ESqKhuhkrjAaFwmvS
MEpEN32p+HtjYVLmVSL1CrJdvDKfDWUo75gSVe1903IaZY/0voO4+3KZ827tPILc2EZuL7kd1ppN
4X7bdqvtx0f9Zzf7Wvv0B0pGKspSL27KFgI3+mMTqyHDhIqHhhM0GhNWNDlkpi+4GgilNE3edwUe
Q2c1RjQn4vIAMRilMG324+ICd1TwxSbwQ8p9lJlbLcxx/mjtDdsJUM0/rR+spyCDYSYFD7XOddCc
LQf4l665Q8SobfRufcMKI3P3iSXDVWST95sZNU63DiXzouyRmuNb2ahgiKiAL0mblhTBTpppERpr
ZOal+qcSWULFN1zFIwNIY5xQC/pYMQM2Q/qjwk3vyacRQWd/QGB0du0+SVjUGTRduJljSwksA9Qo
bjbCwU/tw8J9FkGCL2rrsQKHvYhCWmlBmMrHrQ2Gt3awYfRUmwtGbtxj8weln9/Z9BoTbG/aYPcQ
4moJh+Ma/jKKdYusl/RLPNkASnViEfG7ropzJL6hPyvd5LdH0ITLI4DEuEJkry+5XmEbc6wtB4Xr
dmIlItMY+TOALGkkBCyqlYGOJdS+GDH/uccfmVsBVvOamUD7QJ5JpURINAW/1ECydDlpeVYX+w82
lbZmE3tnwQ4JxhFZHdqIncUk6u0819uGK8ECBYYFyYh03VxWt9SB4RzqEEZL8Y2GRwsVasIpMkEx
Nq/3aaYtkHKEd0aYudYWAAAeKZNrrVPwia4Mi5Jxh3rE+kVv3aAOYccIIbvHxDvG3hLkwxMzpAbj
8bkOShS+2UtZUF9Yj5G0feazz6cH1b9a+28C5mFnNR/j3Nk50j6z3/KQ7X2BgS46hjB7a6GAmgfX
UicNPnZ5UbwI3LKJsyxsQq33grUnfTha2WoftaNaBTz7zZtVHS/apSb7CjSxmfnCmZAsf8qavxeT
U4T40CRsmbtfTKbj2Jwd/kvgxT3VeFusnzdplUTt0rBMeTLb4EDKoI8moyi9oLqPXQCdEY1lWBH0
W83PRcjeJ1fl+27zCo48GaARBlLWUNsVgM2eghRXYvX6RwdPOEzCaGcGlxS9IcVOOAWYWWL57XrC
s+FGE7kDdHD67BpNtGObWYYnXSLqJqMkMWjgmH6K87u93tRyPN2QMO0o0Q9Sq+VFd9/DSOlS/0B8
29njIZh41AHzm1tg7GVtmf9oE15ZAq928Yfdn+AD2pK0zOIP8kEtYJt6tJ0BhUK66a5VfkWku4zo
b3eV1HpgM/qUQ0+kJUjniMB8aO2SnEDDOcB0M0Tfafu8scQhGlUs/BAvsx9k0HhAeTuL49tnmrVn
oRIO54Zz0nFmRrDvR+N3PGhPEogXZZM9WMfS96i6c3y+VidP/BRf583XzQsnapMbVrrTf/5Akt5P
oSxj2awDJoM3kwFoJc/y3bIDnsdDGeSa9osgisd6M0UhpujJKAl1x8X653FNrjH6zj1KeyT5xt1l
bVUKlfb3w3wpNIoZR4C3hwJMWgw0A2s3urc9S0KNhmcZpf6+QAO3G2PQZECR1utSRmb/NgyIqiOO
S1wZgRzBvjeVu9Z6oEl1g1mBx/7n5j8upE1PwSv/5FcbyhwLJwlChm+wQ3AEvhtp9umwrgdGRZD+
iFt0tZf/Rl6OfjRA7hmz+7RrHiCyym381qja0AlcN3k+k4r5dPMRTtao49klPfSa/J5N3LGOrh6+
y2TAoKpCh0zlwf3SuPvfcIFrNYIOJwx8nTJxaDKyQo0h/IYbZQaHe7esNfeY8/Zq4KxXTSvCIcPN
1X1mJQqh3nIB5+W6xFHOwE7a8YqdXZQVBg7m1QPl501jy9Lo4iIfEeaJBnwQqPwwBxF7/DYxavFT
QRxCLXAzQf/7aSbGDpFXHkW7kVxk2/ZUkzOyl2yksjz889wPb37afN8lHifR0nA9SSXp5GzKRUn3
SLbIuENpb0thykK83s9Z/yOl8ekZkjRGno+gfN24WNyrq++EjjMTvZjpqBxzmei/OEVerXNnyNCK
Cep2K+w7Q94sYyP5izuGjJYU8aZv/zTfsIx/dBEikbRhQZXwz2iwRRNHlYTZKuqiyb9WdFhHAUyw
ZscFxKezMerlE0cKToO5EaEvYs0qRCDbPARqKdL6QGxdi4ueMJGpXx86gwKwHU2z2f4yAJ1Y5lqN
YBzMFxnmuxea0q+b/MyQfvG3VU2SOW2X9dRP8ViKYiowo2wcPuy+DphGkFnrEDcpnoTS1SIVSZTH
l8dTSEl5iJGbmv6rCuFYKTf7UTptasWL42kQAlHycK7FIHWch1uKLgxdZkWhhY1ZA8Fjjj0kAEnW
AY08hKtsLUPR4dtLyZ0qsRfL5/mH2uUSTy+ryQd/jTv7WAPEoWlxEQoyeThkTsTCvFcGLQB5SmTG
goropYU4n2yONYZIankbDHJKtwkNBCmDM7Wr6xVMKSB/7X2b/rKfvN5zAH/0T0y10+xgY1qhfkfT
2ux0/mD21jpAyKut+ZlMa2ACBwtIPLBSVknesk7LXoYFCiC+i08+HPVSbKLek7lUUo06osQQd8EC
uGyOctq6RM2bha0lJIhN7q+koownABFfIsJaDpzZOkPmu5BT6vfnwVWbK6j46w1Qep1eiAJyYgE6
L1OpuqfN6mXEOSh4vj5rXOYvsbjkDCojzAp/SQJOfH0KccAglCFqfrvr/888ZcemmBC5cIuy0Koo
0B5pJKpVTlxme2KoeqAqH80vl6cDEmNm5B9cDiHzTvKTMGVGrBItXroZA1zuOIO5UDpyPnExjIat
Xvi3X6AKJlZPsTzLTaPPn1bAp9FzkzU68dUp1mQTeDN5RXWdSRuz2FQAU7BbvccbyQ7DD5NqZUhu
V+zLIgNWqx95JSNxhQvire3YPfFOc9heyDZSAS+drPzoqQndUTjmIENzYYhZgzhWt9Bm0uUP2v7p
GSir2W6ItB1iulI6TtbaVEWGwMiZKlcr19XnZmo8XmTG1meNC9PsVr4dxt00HByQaF+HmddDbu46
N8C5vTNC6TNhzsq6vSNEKchWNi2KhOO4ChfdbQWDvgqDgpb79dzKLcV56ZReHRXgUpgFY4N8xxjI
V1nOhaGeDisrpTLhlevd4pW/kl+T/xlN9wEWzTb/uGI2fSKPLBx4hUJbT7Sqmmqg7P2Z0AxR8qfb
TMILHDtAyc2g+WNUlStZGfRebl5G6EkNYKSDaNSfQvDI0xqajx13sXgVGnCLXbB5gnCW1rvEUtRY
D3v9qE+Bs8sJ7hTDBGl40bBzBGVzXl2nuGSCxz8c+xqaNr8kcAfGGWI8QGxM5locdNcq5Y/jAq5C
VANfX1HyLpO8tErh0yyQ8eUbpKv6osfRoTeo/SnBHPqJT4/1Gs6hz1+NKxyftmqqlePHenKfOIoE
YQcYsyKTzj96pqHLGxfoeEE9KNvBcm4ky745SRCPiyo7eb++LFq+41DDGRhPq7kgiCpcpV2//wTR
0xr98fb+zB6WJWO+I0SKvaL2lcaCdqqTe4MICRVh8vYM5rumaHuV/PB5wkB/FCHB71THti9dG2v2
eNcOMpjMFcb0jNPJi69s0mdelKPrU7IKdqNt0o2W2iClr/fQkrnng79KtYtI75ULaNvpemmygtSd
Z7w6j3S1yGb0wFhTB9usvoNIswYCEJ/qcOPLuRgBlMwnujFczLrAMDH+GpOGqsbsJ643tBwpCtge
NRRBEueet+0/qV+SyGyxXCQC/MFOF2CeECXjOuZrFK6j5MiFXIrsl1v6HHHd2CuUU2TYzmHiew4T
eMQbTv4/1md5lHQsu3AiLHI1puVEpVAqDhflkrIJE6Lq72QSXHl7lHFAL4GLYWOL9chbV3tndZDu
3OL/GOpy73HYqqGUh4xnGkm6B7mIvKndb+BjKZWRAr0dT35C6VswOOuFjHiY2o7d7J0Rl+LQQQi7
rRXDhzb1airIqIYcR861WGC/uQC6QD8CE7EP/tmj/wrz5LXUbXqR8SHgy+yNmNlOR05gcI9hymoI
7raW8xsZJSs98oNzUEYZeqPthYY3MqO6/SlL/y3/C3Tz75XPfjTUZde940DAL7RLiUboHDsyiYMt
cucgzZ2RS/4JFR0X1EubnlW6kk+iVvYPexKIi3rvod5tYj3s+IJiNzqBrmfh9JVezP4W78Hnm2EP
lX92bU2/2CK37aAGQiQivA9RE2bXMO4Nsw73cD3MkhslLgRzYTUKseVndruT5vjKJuX8aGQ9s57O
IJm6Bf1PEBNVODhkV2DDduvQ42Y4+N9QXMMbGGAMaJUBmvpObIbMHlYW3dNPkkQz4ZFuhPli/Sv7
tr3RMxzK2UXCaRiz28cM2Q4jAX8an55kL3l6EYU23nlGj1N0U9Kie1duVWirtdsLIy3ztpEU7RnO
6EYPVGdgwMkFeEhwvoIrKSfW3rb4yRZ2JWN6gGTpKZrqNckabXgk4S9P76z4Hx5c1Dus2UFFAyP7
wi80i6uNyHJOIuCJvGqs4jmPwX+f7mB/BAayUUj39HjUIKPjyHf4vtFWCwi/WK0lbJqbZlbs1ywl
d+hrksDIohSPqWO6u8N14Wds31SqNprQn0o1eyUPGMt8a7k1XeM0/Fsyn6g8GhUz3jRAhkjZ/W3A
q+qNmY/donWm+/xnEdcc/ARxjH7aNmy+1kaivLmUb0KZetJSmy6gPBDFCKtz4JQvi7SThmCBHILF
DjtYFSCiqyZXmJtyD/FkLaDPFRUjFSK3XF+rfydPjl49yxhbuwNjZ4rxzU2t85x0sDduMcs+S8CR
9i3shNHWtgA4QVFlV30GnM2bcS6dnWFGDq60uwbdO6ZTBgNW81f+VkqYVjrtTTBtAE6Rwn7Af6JU
zB5TkZfJ9fhjkZH0a6sACop7JzpmgbH+t8gITLhEzVfH8zXkKutgdEdWMY1uo4pd+mYrR8zZZaX+
HbJZtmJg+7x0O871Mz0+ZLsITwAvUMv+AIGOdqMjTZq1e12vWsx5BjaDTW3L+18rvcM/ho0FmWf6
PxrlLvthTTzZvltH+4QYpAYPmP7k8nzPZFx20PSmBNwKJuwoEGGB+zJD1DgSTTYh1S5oVXwwGGOr
NhCLhBoKaVE5TkKZHUA3NgK/gfdHQ5AtavLCWG9mHSG1DB5i6y3sethCiG1u/dHwQjyzoUBwJCj3
PrkjDw9uqlTpCsEprtVmIJA/RhJ3U8NtCX8aFZGngfg+i9AwfouFVkU03MHsfEZ4w49/Qkjozwtd
wtiDu4ubddDAgkqJpEU0fJY7O/yJCyVqxVSqtfKZMo8ufrfcKaiBhkbyWQ0eYoFaHwMv1s3F7H6J
F23q97bY2nd8HIZXteqzBVxz3BDDSDIUO+uTakQtVPEki57zOEjxWQvUyv8R0phRiI7MLvq9Uic1
`protect end_protected
