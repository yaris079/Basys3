`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Sas/3svv+GFK1oRCduCVjo8cTO4WKln2PTQ9QySudiEOBnlgVF0bpFG9K70+dlwox2ef9Jh97Zuc
7f0t5sTi9A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CquWK+KUo3B3V7qe+SbVFguZGjNMbMm884v1v078Tyhe3h36DZsYx/xGA9KQFEntGifUH0YpWvVW
3qDJ99mTFC6AgAQwnmiQb/7h2SILOmHReSv2T/9KYmGWokYF0o+081+bBszX006Kn9iahR0GS/I1
wKJp6rSCTr3OFrJXhm4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TitgIY1JMFElOVw1zGDvwut+ZvA2WY67VPWM7Ok+Nr+megJPCxt0UpaRvRotqxP696ocRx880Na8
mTzmTgOWVVa8aOoUfss/roal8VBz+DpL9cQ4W7L6e0hX9pDUN5JMGl3dd47M/24q3NKmaoYxW6sV
sIXoI9NNE24MwblkxQSXvT5dyyW6KNPQTcwoVvA+jsOEs8OuQiV1cyoktVVJeTHMmgGcOzV01nbO
4VMUcp7d1N1FGYfRpRTnEIFap/rNj252vQDkTo29vbTrS3fFtCsuYs4X4XMKPfS8FMEeHb+JHraw
jljacodITezgWknhTkpT+iKm5Tqoa0dCMYxbVw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Xmcv/yOMXBA8vnDXw7Nq74CpSXVBIsGTuqUwWtJ+jh4RcyMv1r+GtG3wbI8JGus1ItwTS8L776ES
VQmjupyqVQ8f9FLXXLdD3azKBx1g68hlMU45ZpHIUGJBRjaXsa3oWYNbnpR5ABGUe3n5AoRGz8/X
WFbxNx1lmeyr+Wn/DII=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
oBH5ek051LI0D/v70NPwLobmQBNiM7a83U7zw5QlQpVB6jjNj/jD+/HGJ6/k2FyYjssEKIQg39vS
qwMSwmSQ1QHXSw6/oQ83yO3zkzhgmbN0Jf6BuHrdzdtO0KMqPyTLKFpMtQLTZB9yJCYqTG3r9wCt
HB6KdmjGm9RBM++fy8KvIPspK6k0TXUE6M8I7W1Z3qHNU7SA5qKOLB2/02CFr+Oua1eII3DM3n8j
fMv++ytpQhcXoFiEibSImy9aJcJiTERftXaP69qqxpZE+K/97LotwnD69N8BaQI4Uy//4xsmXIST
lo2/DyaEFR+U7xbM8vOINL5dAa2u/QgjQCGgsA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 54544)
`protect data_block
dbhPMogRuqcd93PeOXUANNrTbsX+btebeQPsKGVWvnZSq16KmF85AoPwiFdgag8bliIsVwIMAbNj
C/SGsn6jMpiH7tVOpMPbJYU4zIb5qZvaY+Zcy5eQSrznlpEj7F3/6Gbvvemk/PMkK8nN9qFSN7fb
KjK5UHHqQ7lypQl5SvPjK1NJI9on6KKqlBlWC5AlZDrHnJPfMtea7u+0OFSl9R3Tg6zS6Q7JakXO
573bONwT3+DAFqYy6vdzK48W71kZWhOCbAac1B7dJ4JzKe8/BAspnrZPP4YpUJABuiCPyBz/twz4
ZSKZ+mnl3OjouVNP9yiUz0pR71+pVP1wCtJyh97TpdX4u24VIRcWjReaUTT/D2wpTcp0W/xXcoN8
cpC1fIBQ9nDMRPCiskVaRg/+LcRTZz6ozKumLViexM0ijA1e/YbOO3rUJYv97ho5y70G3w8XyCO3
4ZS/9bUHzYRoZbZK7IIAF2JQHPJBiLzi5AvTmm7PV1SBdi5WD1aUXwQrN6bB5xKlKsX6emA0eyjP
G8UFiVwqoyMFS5N08/q7cI3EztxuvkSr8prMi7IICWE60mDyXYdYW5EHovf6nLQLLDHvjknXmrku
py6/wtV5IvCic4f2uZWhk1WIlJFeuPsGoixBXA/1sY8OsUG1uOvaXkN0+Zt6cxQbxGiHBrykIdTu
jKhJkuVXSmEru2Zdc6wRtU1bCfJGBTMeOdKu4MjAnsz8n/g4LX1QSNIvqxJXbv1y8RmGiTfApdQt
ksTATYWLUxj7xkAaxrnD4Eh/bjllZ2HmXuCWp05GI7dyi+E+NEvVNkeZkFGziBCI0j6rpHd5Uo8k
bpnFGHRVjbhW9K4E24e/9gP+KNEm8QTv6/OiIRiV1wxc37K6fPI9WQ0BYS3g+rnl+fcfJ0T9RpFR
cdKqntk3ns+pb5E2YtUi3PTbKvxWAuuOL4qHbBFFfElX5N4PD040xtcLQzpDolhIMWDd78NIrprp
ve0blLl5S8XPBK4UCP1RN4iGWurNSwXPIfwS+VzhGYopHuh8Qh8mreCp5Rgvd6cuRQYdSTR0M0VT
YRIufTTFtQVbeSo/oPwh3pGxbIfcLLyeQfMJ00EKrLkEZ3x/t8flpr9z5xh9MPmFIckxhbLN+a7N
fVXH0r2o7h98V4W0gmQ9SLPhQXVzEF6riM3Bnxv/QHAC9tD2bYcWBAgERaAWNdVJap9nMimjx8cG
Qr7ZjTh6uEDYCD3n2vB4DapXwgx7cQXTCx1WdrbHCf5xiHoL1TXrDtfz06vshf9sJou+bFY1BBjR
yy447wRt/pY/j28TMWWdTf7MrCa4jrYdkt0vMFX938CGTP5PNpCYcfxRI2KrJGo9CmFyysNextF/
wMEAsMtiAenUA3RnbEP6ldQb7VPy5+yq9C71G9GFGg4Pvqv7qlM72MVwOB3Ie/7mGuSZ1pEHTxOC
Bi9IdCYom892pfJb9mIGmXSo2+LOTpVdiH5g9/p3cInWlgGu1Y+EFoI9wrsBA++MY2Lh83g/h09e
4ceLhX9SuoH0sE65fQWDKhfbgbLMygaXilVRd03VJgPf8LCmc6IBWyDM3MV1VCOT0C5j705Cj9GL
9YFoX5xKDCYGMuG+sZXCDsY6ZYn5n9+1NvNVjnmHqRyJEkLn8yMvifnUDFKs22MPm0km1JOWptWL
PkyPt8hvpVgW1TU2WtGnkuJaWUIIazA4smMvzbWuRBlRLOj0gwN8y9w4jLOZezFTRk7atjiehq3O
X+ziTI45NYdEpEoudn5RdAu9bptAOgm+vQgzAN7kdqGdmRtgdEQ0d4raOpg2GbmpL3u/gkNRhtMd
4DJZFppiPWDNjLXDHYxuBBMah1bLjdWFED2izWl+YmLPQK2nANIZt92JxUVy33RffsuThnIGRR9Q
2iSIncQPLaqeY5qMs7h+ktHQsq7IY5c1Z+TGH8M551YEyQP65RLq5lxurDkXbW7McyOTZmi25NmF
rTaHCENDqXU2CWWszdoC7TiWTmWUKcBY/Pbz0RNBiUmlw/B175vemqRwntyjKSbVDeG125iNi5QC
i/Ot5sTVyuGEkqXCql7uomlkLBoVRp/g5G97P5YkUW0lYf9noX/tjTlpnJDBRx33n03mY8tRfGQn
Ku9NTYNudFjun03/+sEbHHJW29jClwkcFqAexWvqW19UD6Jwf+/TX6q23R/m9lRdWEfUHlSXvafL
jQ60yV4/ONjTv7sDUfT4+5rMpsQ+CMehgrMzxmjDXrEr0jEhRTIM7XdXr8jcQjYJmJpvGmUoMetg
srySba6zgqPbRn2VmYakT2ccB9CycI/DjC6pKHrtzlVlmHPPRDIetHLuNxN31W55gGgEwHys53Gm
EfrAgxtgtQzGM1DAj//aaRsvdza8+otHDXOz9Cl7QtthRmzvekowAFamrqousE+YlgidKIwIepZb
b1ofDwsSi1Co811HFoIZ55lopfXTcYt9k0GenF3MBGGnF3SCl+So/WxL0Jm5Ienrk2hGFBwLTkYm
VEGP0kk3CbG7F22c89dNxv6nbJt9kUt6dcA35buWb0DBzVchPl0YoeQPbjlmL7YXqNVjbJ0nAP0a
w8RjLY8MPvmIutqQMSRVRKKjUzEl9bFH4ZNEDtEMCK4/3oHqm2xGyHIpcFHq4zalmkmK4D49gB7G
R0nhUSm8JoLBuf5q/BeoOYdHl7yD+9SPUKvyxFx4P8G7vge+C+jEpMkSdEviqu87/gRpavrZ+H6p
eoiRdo1Wn+fbyiHkhL0JqKMlqrsxhikVRUk0v6vRrgRJIki1IxA3Y9BR/PlnTgTA3aRucAG6DNvc
qBXePvtFYXmiOLbSeo52LnnGbu9eJtqSL5zUywfz4oCVPLO4L87GTAVSrNc+hCLcpNYTjnWu1Qag
3cxKCKBotj5gp/1IlnEhmoohoo56ubXH8S/dkab55vhjK6rKSSInPMquIT8dpm1wVOEt1FI6gE8j
ILrfD/TWUfn8ruhSzFiXW0Vye+kkD3FdTrBCgRzFbrLsolUFfig2cJ/jziY5mvUVWZ303DyJu0nf
zs6XCLTVQ1hS8M7twFNEGfFrmtB7DbZA1GWYuIuB8r6u+o+EWqq3aJ3Lezxy7OyILyoJ2zp6uCew
ZY5jGlBoDUv7iHxMLz2Uz9hEXCvGdBmbhkPgmvEI3EvKGRNZTs2kxIxRLJ8cDPD9r78GvepI3PzU
KvAQltEqcW6SACEz1IA5NhWNzOs6gdUpspFrb+WNODceHNIBsWz8yIwQBmu+Fs5uUauVZnYcF7eY
hx8o7uYj3m6ZBlNue6mlFNY07S9nqm08fPx4x7jvhkWvsx7Khz+YeyZsow9db+ISPoA5VAn1V+tF
G6+bzYo8D+fgv2CjpLDdFiXOtth3VBDxdNlbF2bqWsO4syGVMaAwWijQ4XkZd8XecUOxntssYj07
G0Nbd4OWaB2HRT0qIcvFfeLLhAo73/p7ghMNQbWoxfDZ85NvlhMB1QeZI3V7Y3IbpJBkngAyC0l4
Lj1feWU+nIDO3QRg7N7LLFfLJ38vhDgiqmtfhMydS4tV9pmiX1xZp5JToIPRXc2YcW91vfwDbjpc
UsFrh1mfguQdLxSK4QkBRhCPIljgHlGL7gKx49VEkvP6aM74QKcbyNKGaBrFrzkSb44W7AL14TVm
BS1v5QyEIJRiUFa5QqkjIE896KzNWnpmnmZN/t1RAE6LATQ3ZX3+7Wt3JA/Jx5y60AtLkrqjoABP
KhN+eEeCr3mqr4c4ac8Vr0PlC5Yxk/nJwfubclngzIka/oNKECv0cXF46ReUvqcXC8WiPssFf7Ha
5jRZF/hfvMDUYJKxhJ3Rp4Cyc9T5zNMv4h3lO/5S0ZgLmCfnS8WrS8WoAfjMLR2bDhohkLUIKxgA
wKf7iaZybEmmu6qYfR3n9OFIvz9LJTFO53KpFYSGYRrk+3/vMco46ujcSfUXTwLnL79W69r3QEB+
0U8Rm0W1+Y3Hmc0Ud3/tR80sxuZONmxnpNyYazqb/i0+o4U9ngsqsNG4pxGS9k+BZTRKu6tQxY4N
2YP1Ly/UO7loz6ysuQwz7mX3i5nk77Aj1jHXnbeo1j1Qafi4O4wYZ1L+FBFX9tziWx0tWYYuVp3H
95o9Y5iGDzaAslq/BfPhrzMZPgMxHCbonkQEK2Jr5PDv1gcFuIm66bXIrPf/nrlDAtUo4di9hnci
PpOWSOSjmIWbSLgKT0yCWnktKhRPeraXlZLyia9UNEfcegCS+ojqu28BCEROLhBUb95o4EJY2wrl
oF7Im+ubfVORSkq8QJVT7w2CHFhgaVtDagBIQd/khRsO42zarnJ2totkGwZKGaLtf5wZC/cIzF9n
/nIzyeIw1rGXeAWJ2iwbjxEVzvT0AqSEwRlEiAvcndrZN0QcmUy7UUJRPILaISSaM5ECtfgnUgGH
RpB4XL3rircqCkFprujHfCnrsXndbk5soN4Ze9E+/PKCiIIpjdS4NWDFpYpdxLpTeXEaCdI8MaQQ
J27C8wpf1s8YZVcRjNjZQlqBgH9Oe30AVrXdvCGRGKJG7Lfp3QWxNjJeHQFvD1P+XMJjhKhyQR/w
Yp48K+jeVuF0SQ0uCYTtJktafGVFlEDYvh9x32voXntz6ruS2ZRAWPIZkOEWsYT2yCZ1RjmJ7ixT
DoLoSqNKD/SVBNzsYAkspoYffMJsYTNgzeoGEDmimmXInTHYr2XAq4Hl6fbvAvt837ZDGN1aHewI
1E9auL0G1Qgq1UX/UslOlTKewV676OoaFTgVvabGZkBtC8A1CUO6L2PS6jZkuQ8sQ5tkK+BkSHf9
ExTSlplfTmiX1q9ekQGlcbjnlNX0oM+lLfJ6INXT1/cMryLa6kUfXo5u1f0JCIe/FbjfdNxE4zso
P1k1sT/LPitaaC5s6Kpqmobc82MtC1MEQYyL6JlS4xZ47XhKiAM3bQxf09ecsCHcSGtdAaEIVgG/
BAy8/M6lSIaHvE+eyfrXg3TsXIJdnHWBB89qK2cBv5veaWhNzGKNOnPpuLLL+3AWGJ+QOZi2hDYX
GE2YCwzsQvc6KwFZsv/4nYAGAjiRVbji488kkvfrY2DJc4AwZn/JM9s/wC3DRpYDJcu4PrVnFiPE
SGw7ndt0SJadtaHKi6KCTh2BQIhwAf/IDBv84V3joxpXnRj35uc067T9Lh2wz1TRWnSPJRM78IE6
VyEEXblX3wRu+svhQCH0yhJuoHzT4aPRFT2jX+opDf8oQjvfJ/f3UHzDu1gM1UL25AEpgpuCbRQl
xtG6YnOlEvkybbfDeYuXdqM4zrZ7EkUyswBL+4gTj3+xQ3EefUu9oBfNQ86KLJsnY+ALHk96Viic
StgdQSl7F61DSX55K2dQQcjZCYPwmjMVwQINTx2Awm5sxE9cbVHMWRnqSypUsS0plmH3keBk+K+5
C9zweQUQ88EqYMvBLYkKxS/fRWxGYgB00g6fbLBkJKpNjqSWwCsO7yQGTTigLSDyoiPkeVrnaegz
658rFvcyBli3tIbo261/r1h9uQVK5KSeWaKIqcbxn5VLDSb8VDQkeIeFcY8HgbI4VAdZNm7613a5
bJivuAtG4xiaf3XnX2Dihe6lP97jjtnFc1p4uffiF5FtyCpn3GIyCwFNvO1MfhMCF5CiRaDierNE
gHjlEwE0N9iIYkkrGpEIDx28SZnCgnCfiLIoPbRpqSo48PbedQhRUMjpYSVKVvFyri3TWFn9Lj61
zXxzpPyX6xl4Jbb9vfUcXglI1tz6uE/JHSXqrtpoZVkHckATrQxMTERuWXFLeUUM4dC4BIJXC+4D
gD3hm7nyqXLB8DLjK0CyBTwg4FJjr71CWjCglORacSPSs+mSFJFV090Cy+M45+12vq25ABM6mSD4
3RNgjQUlTsK51/xvzUKmsXP/DWYH91xHCh/eXa2MHkgJLP9zxiMJQ6Zyo86f7Uc2JflVwirSUz15
4BHM97wYywQsZEgpTUCBDMBySpxDyHp5DLaJYGGyCTZT3pQ3I0F2cH48jItXAUXJlHa1y3SaWlQx
QhRAmTnzww0SsIJ86nUhMMfJECjHSJGgR3GkGxKIxDM638I2l9VDScs7lEOvaHRd19tAb2DY2qrD
fGHm8N647P9Ro7AAheoGQq0evjgkKTzC7+DYNUY8fbfijFZJ8YJLdDU9ehNyeV3o0lQxuzc1Ez0e
8sFXS7HPogjG5NWf4R2txWCc4RpklNb/wRJOagRrJqEjt7UPvCVrK+w6z1QunRvzam+gmoTkZlbU
KvrH7MGtwTFzvKelXNXuXtzwsoLnGN8W0wLhRY0tyqWrormaIVZegTQfPqMhCrmryPAgV/Zt8PLh
TQiUGJrziKSyeUxPX/Q8YUvr6jeq+6Pzpt21vJdtLgb3pp/ik1gfXHlqskIIjOK3iDGufjHil1cA
9lmug4Pmn5p/RFS2Un70ONzRsmm92J5+E4cbwUww7+/yFwDMv37ULWZS/5DFuZIF+tOgHEO7OSLk
Rsy/8Uwon7kokKkilLUYnrYXMNCOjixVh8rYa86QPPO0ET5LGFX++y6bpQkNCaxqHpu3xn0xOtOP
FDkF2R9tuqGyE/3o7PYoZjb9bjWGp8ZQeqZDid+t3YxgZoDDhP80ezvm8iV6xxxP2ozODPsyqC+3
hr4KeUelUZPqvDfyuu8a3GRJf6itfk4MlWEnlMAZK7FYjwc9No0/8BJQ10aJ9ZEKExPeZInd501Q
/MMvF3C58y3GDXfL5H0MTqlbzWQ1bKa4iZjnjjMKkJjp47DMV3IdAf1OTDdqt0kwpSyqlmD13XWZ
M9434MQRzSQaICcacD/BgWd9whMnT6J5Wbcrwsb0JH19Byw7Lp7fKZaD1qPovvjP9eDFiPJGotWn
GnOnymboqsMOccIuyeairRszAcqsjz6r2hwzAuyQjLVUpQ9xcdpsWtaqx3QdnC/hOVqLLQAeJ/Rm
EYT7xHNz3KLkz+Hy2mvtT3HznP0MiOLkuMFGyemH2evy2ilLemBPML2tPdoNyNc4X5drneSphr1j
E4hLzM8qwExIrnDgLPWZ3/Ty8slKskkkf5cRs9CVndwi7s1AHsU7XOyKwSTYlfROB/a+9ug/9aqz
BxVaeBxmR78rIpf6KmEIbXZdMrFsj0q++Zb24ktTBoyvC7Yzoi1IaGX4BZAIXJ55RtJAzFrnYaKT
MIk0S8TJ+EsfHZ8xDMVV2671bC5Jq0SDDmAUg05BNVnjfATMU8xfgYe47BuYqdyqxzGXUwqkyeDG
B/5a1dVqaFC0edD8L3V6FyU5gBSNTxGN+CE7YhW8kG8rlPPomzpc8N9o5ob+BlKkHShWsO5Tt43n
ArSbKdDN17bKmmIpiA8QqmZ94X/57/kjCmDC3zqbWMyccPdyGWpgBU88J7z3iTlkhKcyH+ZtDijj
Ge+gxsZxu6m78HYNbM0PC92zUvGXYsU4XofbhB8U2kbcwLjy9ZOkNq6GYRkm4DsCj1ue26F46yMI
o2uTctaBanDuJqCGvk+ooy8PDvBKVXQDvJurnhHaPDCy0d3B7ggZS/JMK4yaJKfDeu94ULHcyhNE
Lnm0+fCqrkCdzayy4G4RYjDFapcfxInfnhj8dYUY05wWajBGarV2A142okLwRKDhiOX6eSghcNJp
HYh553CJLLvMUn0mZo+Z0PMes7A56chRRmQeKJ0IiBB4xrcVSqu6nzTQL4Eivi7YYJ7816BGpVhn
TZLwx4I97c/OYSDfvIlwSL565EYTgVlpvdEQQQeltORwqjtgZ6P95RT0Q6cuI8hgskHzxeNbFOEq
YfDPqDJdSRnur+Cmq7rcXb7ywM2itQpf0+gMfErBZLBrkq4W4oEC7xIdEocbSvK+KNckQk5eoZUP
3RnK2BlO5iQunMD6rdmFK9mMLodX/bMQMZ6yhSeUvvkGISex5AvH6JdWgcRVn4u3clb1cXWMTBRe
JkOaK//nokgp4T+C8eA/aX8OOLS6zoAE8R63h6QFSzx2d7VP8n/44EmCgAXE6hqERIlBAeJI2j6f
w+iXFDP5NKdBrpQbSgXMQZiB7ZbBwtjMCB8/xrVDa4YGJa1SJA5dZVczRRhXxQCOLUuSbD/MFF3q
tsvgJ0tIc1Y0c0/RuC8LXY484ERyn7LhYzDCWbBBZeyMB7wUNfDAqiyl76DYkGTw0HM3kk+mpG62
ZIgnucVWslJDNKR/k2U97stTesCCiwFxAi/xErEAr3q52P6ELczMcyqDlzWtWD1vOfQkA0ew+Ki+
85DsJzbv4Qcrl/+Kyjrh9OxYQWfp3ccGvhF4cmXtYZ1iEjNhWe3OloHvOWMl0AyDKMljQpmHcNpr
CNLmTsvI2OQkUVgl4Yuuyp5HK9bSH/8+nQLj4ug1kB8FjcNkLztLeOvsrIiYWecATL4wdoTwcPFM
S+IoONxnSco/aywPgiYPE3/fE+QbB3JrUFPB0jT6KWzQ+a3EQJcv4l8bLlBvbalBuCACeevjNfsJ
uQINN2R/oRF7djotrsTss6knXaJix4/sPCG9cbMahO9ltuNhf0KAdPywF3OfsRG4kb60ZxNd0Sfq
QpgRlYIYxILXsmBYjTnAO2yKdtTQJgMDtbMK1EDliSO9gaK3p9v5zQs2xGUrvrvy+abUCa4pUCeA
hrn+MEJpbH6WhpOlCjJ6yODz0FC1w2O/AnbRWc1wFlNeYk8Dp6ITm6MG9t+PvmCiMEMUhz7FqMIO
aHBit2PUp/sLGK4H3/NI3G8ziAhHTt2A1c1wJ3a81k9Oo264J2bsLpngTl0wBf45PnjS6LclWYRs
+bcCauaIvzvfAdLGUzcMEmUJRtpkuhdxesegRrSVhXy5sKHuKujsOFJpdrYa1+B3vVY/nKTtHObG
z78UO1Q4pS4eMSXaXf/FV4kvQpwCEO0BfDzke02J6jji0bpqn6kYideImYqHuh/jJWhVqmlj07ed
McbXlZZcDRrD5YAK3uj/ikVdvOc0U4TOgKp9QDA/56o3Ve6eWykuQwv2BQsJupIkdUJE//hM9vIA
jK2Mi4iiYzMIA9/uwR8Q8t4eIHC+S0h9HGrT7Rh8tscX+r84sOcHG9Tk1j3Q/x6mKEZRaMtySi/5
YFaM5CeyQ7gkA8c/dujyTWHGaCo0MrAM89AxLEysMN8HUwKXyHcnwnqrT1P+djj8hgjM49m4Mv2g
Fmu+skzUYCsrUW/atVMILLcuOWXjdRYjwPUCvtlV7dMvd/dcsnO5MxquaFD8Rj7zLvgUp9mZ33zy
qL/xl0M7b6gZ4nDWut0qucSP925kA+Ii65IJ9nKwzRcMbQoCTXX5N7KWbiNAZDct+KBr7G0jrClI
NidpD2w3/0aKi1Gtz6jimvw73wyAWkyk3MAazjp/LZtczPyIq00yudZU950X7S0syylwPErSaoZ+
1H8MW9feWSMttNgTpkoeXqyOudmSZXmsq8MFdrUOVc7wG8YJ61AZiW7l3OUdFNc9lGehWj6K9iIB
LfQ3gXfjcJMT7D7TskDmdEIeFPXEaDz+u5brkTRKftykLpTkufufNA2Y0R9GWU5ZboFNM0+N537Z
G7FFKvTcUDgBgN/HwlKT4dsEGcPkBNhTAARgE0loKzFMSzmP7VdJklNY6fJa0HUlJhlIp0vHxYnH
mhuorHj7KwsbVcIrvt5AyhVaW6b77mxd5jDUKanywW6mXH3xRV/mQw5IOUBtSF484Z6V5ImDiRt1
dsn6zk+6CUTjXxZ1XH+Cc6/UIQoHzriIFr61M5unebRDL4qZsXdupCCN/U56SoQ0VN4cMhqnwYJy
P1HVOc7wpekP7v4NNm8oC16ApoJdqmHu4Xj/7bJR24d7Qk1n1OjWv9pvX2g6fKzfFU3I+iZDU8XJ
7/Vxu0SawXlxj4bz97Y2kKFQZif7RPIudZGUyfotkaHw2+H6s/tElwzi1Te3YhNJH2lhbYkZgZXV
lleCIipBBRh7zOXvt1Kg6YduXvg5GLAVtjnXWNMueM+OyIWgA4tygBL2gJznrpUgkOC2lJufYhdZ
eImja/95PxKEb76BqpDHOQHmGCk4UasA7xJLwUZUT1+rgeFR9vmgy1h/hf16D1BWg2dr4ZrWa++b
8UAIEOWmb8fslbEjkdyWx9K2QC8RLtF4pCgaGbmz699WcgDFHREfOhGXDmEVy35LJIP43gtny+wm
Omg8h830qrC5hwp21Ux+VDJN7IgqCivRqVwFrspQpPUzWk/ZdlEdrtK1TSQBCyz/kMYNW51pf8BH
/4VA0kmEWY1HGndY4c7nwMeLVhGsLMkolOHdU9Wb64CW1IzdPzBd3Qi2W+huysAzDq0RiMXq1uXd
U3CKUy8t/TmdIX0cM86u4WVC4FZVucFOP2jl99HImHYWGIOnjUR2ofBpzoMqpfifqmMPpXcsiGTG
7lyrP+/hm019YbTarOhlW2qaMPEWxY34dYB9atGsx2LSErLYLCVVl+mwjYJ6f2/Pe+JWk1S71rme
LfSQB9LiWtXLV+MAGZyEJHCeR10Euxr1nSiaM3thGnYNZtbd/v8+iCZ9hnH59/iXk22xMBFM171b
L3KrAgKJXlcl4+IaDTfW3ZycBMV522OxK/Hj8s6ubPDLOYikPvd3vnoOLkbbga5paq/Wavjbb4bq
92cbzi0V0X+Mtr3S5M+ZzeDpjfKcdgZwHTQ+FSpPIlYFdF6dpptOB81SKbOYdgNHXaD3S4IpD2Fq
menTgP/SYq7lMsVSiLR7MPpjVpq2344yTWnnq7pLl0FuRi74759IYz6z8r84UlCP38Jh9RAs2eht
naZuYqLWoKYi2KhhXOK8BlZGvHa21E+qoZzPZ8CRys2x/l3/LMG5MqAFukX0y1qL3SybAGhj+XyM
TAEbv9pzcjTyoQ98Twxzv0iUuY0WbLuIQnPQYY7IMlQLoog8vxtem6ZXFs4kR7giXa3OfcBm7Jur
/Qt7qfm5yKoUx0p1KJJif4FJeP+6hv1PLvA0Snb1N/PbeLexGSRTg6jHFDxhwTbAoswocmTNAy/k
V03gdRKu4zTYmSMSTxo99VQxclkKdCi9sJOxfNEAw+cHAa2n0APFHgyeos0d/RY4rvXOmglnPpD/
17gXw6L3rDTThyl5HECcMKIHEOllF4BA26alh/dZrgPLJI0cm+XdmmNsMbke54iL7l2lcoynywkV
LKQpgdAeS2Kq6+UX3RyotfNG3utWHhpIpCElR9r/f1cGg49LlrggcJHmAWCceqO6cNw1vFWJo7ze
HOsiD4wIHg5EsMEPwY7x084MWfP44gx9mKPIsbvuwRaLxGdWpdJK81d4roac+yhaPgy6UZ42knVp
iph3a5YdTzwnmu+ikljY5QtUmBqua6hy7qyMilVWOgZyAy4xrko/vkW52JbluWyd8xlgaobooGGt
08h7PFbb6DSb6LeH/wrce4PZH5nFzrvgWFMTK0m0y7oGPR+p5uzCpPeE/ZZKcAKo0oYTUb6ToTTC
39uWLAuIcsptUQpCjgl7iiHsvmViqU5Y5B556m0xgLuf7DXJlnh2O7C0BAhv6Wc2CgjrD4kl5nKz
vJFvJ3iaYDODDJ5AuaV12SM1+WsZ4ivJBCU7Icwgklg8vNi/+5pTtkrAVIGj9s7YMQLNqqFVzqXJ
QNoxUvI6qSZ19jN2dWnycJVaEjoS3Wlms9syAG8OrucqQpKO3ZZVpewKFiEVs+37fhe2ErrV+yLE
AkH2YNCbzg0g/XA6Zk8u7KMTy5am/b1FNa06jpWPgp+6jcF4WxKP6AL8pZ31EcZF1uUPigTM4Hu6
fFv4WPqYgOuqDH6e4hb9LZbkp/C7XMZH2VgMPPVlL4BbwZEmSSqOZDV3bLtC1UtnYMx0DM443DOz
ZPUTJungnsGDXNrnQgJWm6hOwxEBgG5u4acSyKSfV+2u62rD4clqdzSthHYUza5OkIY/penxlVa9
wg9GMJgGzs+ilikpGWBS5eTP4qRod2c4Xi5ii2xI5vdR7u4TwQw5GkUVCZw0ovqq3CDAgk5SB4sn
55ZI06JHPKeuks8/ALVEJDA2fQbIGmr9nRr+KsoN6q5wbpxY+WOlimm+nksTZrYJ3ER80o4+Mbxt
Ian30E2vOFFK4WXSPo8JQa+d40CSjn/Zb0B9k6L+BAm67PtMoAnvQouQOos9CxZW6HcNm9jIu/Wo
BgfVG2cFktdjwTRQck92UxGl4rme47D27JyLcSp7ge9cxr1g9MhLZHR23VcuyGT8xdZ1FoBmgBSu
9DJpS9zedcT4zNjixtvkZ3fO9/gtH17BZkqRQcOJACqgfZaf5HW80jOB58RA1CJtAegW/Nr3a/zL
cgwqGCclZaqaWl5riieS02lbf4znU7OXz4f1jNESAN48hyCFMzATUMkf594vEsPtFzk/ZoKcjTh/
TCtdqwwfRleEozypuiPhsg64IeTsRwdXVJv86doCtbDsoJUiTw4DNDgfLAOgmnkhck3hhCPexPvF
SQPKCdoBVlyyf3GMIVgWWZiestewTt+esmNtmh/C0kK2CzUiGfXNLT/ebiYWX8scBgZa786A52OO
Ngpmnk3FnkMsrfwwd63lxrydgvz2i8RY6nsZ/cZkHOVjG91x+eTJdpc69AsJMMx4tg0abb7qCA1L
HxgQI6GGFt7FBY6rucwSyoCVdIyISTh6QenFWExST66HJfDStk99X0/kqt1sQpB69GdqN7a+2Pap
W/ktF6WoQQ8xD10lS7nsfcGEc5awWlYMQ9MhdqJjO23T8gkl2KqIycVCZ4m4tbH4emtLo12diVTl
ZgDHAeaxdBWaEhe+wNQo7gxD2QEBYZq6BxWX61LgVpB4xKdVRiV4rCdyJEmswmD8GFSaz1XB/SJp
NwcNQAw9Fo+lvNWZVTByhKtSqeP4DGYQWsE+lcjGvhz8ttBxkV/lESDGGBGdT6Y6BrL1DZPMPnci
+u7J0UwwQsvZgfBqhzNyyTodlEFpNQD+y9jBfZKKgGxecr+DN/O+GSvgnnGZnW8oHbE5jlA13ErC
78COi5QEujDxp+RzH43ql8IOcw6oYZIzr4Fh2AiV4+PkNnGXU3QRYlXtdbwkrIllS3GGvnTaaydW
WhOX4TrU522GtkcXjCqimevbYHYNVIzAXen8DI/hkru36lrASrqJHPY+0JFmNCMfwvI+9eCb8WGO
dagvclQ4N6hY7Iwm/DNWoVFLLZBcbP22eD49C47upQhZHN4/vfazD9FfnT6gK7BSYzoUprz8Tj/1
HW7YvYIm/jLJ9r4Plz6p+VELzhccyo0/lXxGokpENHr1ybuMDF1zLFv4UEmFUPwOim4dNVyZ6Xsl
KbI/xW4X/EHLanrN8q9oGxC6wUX4U4sivVJ5uc+bJ4SNmfPCC6I7AFfymAX4NsubotnpAp9WMUg1
L18W85eIEgmC0JZEoWC9/xLCPKtpp0BoEFf8o8RNVS2SENUK1dYAEpL4Fx9NioYGiK3bcfrqUcgI
poA8CfqCwNPOPWQK15fofgTdnY4tHtGf3DVYm2aQH4X0jzxf1Wm8JNZx2A/IsBc7HwH97UWJmqnb
3MtbLeOIniSvM4a2XSwMbRi2dlJ3t1lYm6PK0QoJejnToGjgiiH4jTWv0ZAr6ghcTeOZ+TCfwS7p
w4XIc/DfTZ4USKlFloKcPuvbQuHg7HcZhge9hX7v49T8GSIl6gV+pGMehcuA7cibayuCVwXKH6KZ
7YQrsmDnMkxnFimEopG+VBxB7DC4vpp9fMjex4xUHeLQjdwfta2gD2KB7rN9ektiOW+GuFIx7uTy
1HFlG4ZECQDsOGRyyYFtLNjWxHjzIb4ayFUYFCuRMRbqCVv++tvungyD7mGWy46//pCxauoOsjV7
Yh4o+QBi1ELN2zH4MIBSleYmflNAst78zdhdEUJezR6fofqNUERoM8vk9c+Fd+Fo27UDsQFTVIn0
C4bZlhUVT/sQ6s6FLuKv0W9ReaARHInjwUGtwTms3En6tJY2jWrwS35FvlcKmuOoO4sl2FA2RWZ/
pL6PTFydVwtZaKILL5oAgvfY3gWf7QUot5GDziaIdwquFIkh51VBZ6b13Hv57R6AyE60vO5L9La6
Nk56fL9ceoA0ZFY+4gBUAsmNqcxm5JEXgN/jO8/ghiV+h2nsixpJa+LDeuliwOYJyK1/G8hua9yq
eM8CzZnWHLP2MjNc3UnOv+umypnzxgOGOYm2VtzkxCKeeAqcIpFXnd6Kf8sIGnVWc/3iDCPfVeny
hMl6L9kmEKVxGs31zSe3Phk8dtxLE5aeQ44w9tkR3NVnZHpQsCzvwGDXXN6Dl0/5OZH7V9oev4Aq
Z6w2JNar8AtgnEqsaglgZ68j3H5lYqmdbUokxV/8bZ1StDE3AtaMngdHusPsFWHIP30/Ln9KTJ43
zcz6D8sUrJzgQoipu87oYsvpDuq1EINTRXqt/O+Te0VfVgJvWiMRmnzEn4598HstAo1lMSooElD4
a5R0eqc8gFH9xSdn1FQfEBFKvQ+M4waCW5pYFq/w97M9QLyKMBmKGbYAF6528PIno0v1s6+zO9e7
P0qwaVsxWkyB++jaYNqHUp+8h+ZmRvIc+cOD/s9cIZUlwphmiKr6HPfhcS+9dLeFsoIYqYBSA9i1
DcAxv6DG7wdMYoIHqVATC1T6Mpjvmy9JtGRWJLxfbrYtJwwH/y1hFkoOlEtPdRrpwhpAOvDCpGzQ
7X3vd6Wvk9cb/av3+56mPQ3I6RerrnKRsIlYQB90R1Crnd/Gtk89xs4V8e89BWJa+C/yFGESbUU8
7b6rHRLzxWCD4nQhDckM5/KFw5tZJrfide6oYTOBuGAwY8R82eO6ZqFNtaRb37c6eTipN7DDR7tz
8sr3n9Nv0YX2qiz1VeQZiUK8x0MjDYTPLXnsIiUugdshv2ltQpXvbdPEK/+BArSC/ye5Z7Aa/K8O
v4kxQlyTalLzm07oIqAl2IhVdDojN/Dz6gr7Hs/dgjNS5WEQlFbA1juEDE/blsXK6B+xKbtyIGY5
mGuk4H0quZCznzkObnT8LHPv6sEln5dKqZZsDCUi1uXKyScbvHVqMelJQpA/HHYPpQRggiXQr7h7
EE+4fF1a06z9gmkuTQqtss/dOnVmqTTfQE2dmIHp/AsLtCUQHgnCdcJ1b3CkmSXRK3X58j3cSu5z
n+kMxyzyURMjr6UPsFCwx2ECw04DOexJjbS/hIApFpr7UGW9+Fa+ufagyWkmR8GNmNSeemifCU31
FXc6RBcOHBuDq06kRUy1khrDxkPcYjL+wVHZ6aAadlh5rXgmH1xVvFV0hSkb8v/5x5p4rh4PRAZ1
hB+eT9We6qZ4VnETgQm5GnFIa5Bq4j/mRiDZsC+RqJdCKT/ggOtFS2Xjb9DLJlPO3HL7RW2oG+AP
+phFoZoiNw4QSBO+fI+D4tqiGc/fLsMXAUE14taThewArY03uysx98spsln0y7c8MOc6tYgE2ZV+
EnnROJqsMZiAS4HW0JJnp06j1kGYJKo4zrnRiF0PCFQjEjpHrEH7y+8hHpPlizJL7Vl/0gvyXgkm
0ko5Uqn+3x2RYgn72Upd4mCVR08Ern6IigAlXUYHNEPazXsdH23C1Cko/qPncvaYAw5vFFEhePjL
XIt9j1lhpFd+CAe9LtF/5cWvMVPemV2a4bDXR4Tb3nq0LOP9ZSzNmBZAvfCsdgIsGdBYdyNKUhOG
XiA2zyC/a9uabUr5BFtsoEVLQSXihAuAYcTc6pxHFSVEr2vJTApHPJ+aD05eonwRJO3FIWQHmwkB
OgRik2PU73dVvuaKQU1Rgx7sUeuD4x2T+IE+InfXuTeCnxqWMMUqrwONsr4FfxSG556qm2L3Jj3I
bwpmLUy3hhfNli+0kyC1v+KeCktnrhuMOxxijP3sNn2HADVawMo2kQyLuHqruSKiZZ0qh42us1i0
fonEi9p1P9Lmj2ke8rKKMM0ao5Hw5CiHBnq2jxbXy4U0uXHbHAQgBvZ8zgMNJ/Yfvx/oxo0OYdqi
julPDINf+x/9of4YXMzsdsmxsQXNLSUz7fxyCeSUEk2zkR0+SM3s9lm65BMiyH72VKHOwejS87+s
Dch0ZJrWf7qPoDc0xJbRaWP+SNZ5rcDjgE+J6Y0wDo/wyuX9DIO2xYZkagmQfZlNPEqgMCNUx2by
S5bZ4CC063sx/XSlLgCmrO/1wqhAme8zVYe5SYeOVi7DEJ4rJjBULMKC/qgnumCIeCdu+dkE9GOb
P2Kc6XgEyjfYJmT24h5gQzpI15DtTbU4fzX1dIlazD8TkKru/gq9quMqMszbVN8UjSnefjr6rtrA
aO+q1hGz9uE1NnQtxMR6U2P8flK2EYPEPcLYP/wSIyU9BQrDa4Q501sBmx6MwXpl7+vuoxUBDKaQ
hnTXtHRoJM6Li+gHYtRTNlNH1F85thAiaqQECKhbc7cteifzewk6vf8/LJtfoMgSSuWiRtg/71E/
c0UOH0RkC7rak5BixYaN5RdgUxdsfp/yAC94rtsVruIB7pVGeNdHpRWTq3SBaLZz5HwSjJj3stWe
kjm22O3ecbX8C/yUiwh6jEJjY53vGZBa+5n7jgmpLzXP97VWh4eVwVOxVyvQVETARm+N3XoIyKWz
b3FQTvNBKpTgff3H70/E2UUHdXgoU1AVt/1wxGURUfq4RHLbNnHOYRWRvCqW+kcS/SJuOd32t41R
cxXCqlnMvaTc7bmHGp7Hv2WYzU6wSQM/pTkYMgFK7DfLqbq6gn715ayeFvHOF6jDEradrOsANGCp
co/CNvcJ31f1ixBF7loSxsVg5v9qEqMqLCvbDc9QIImK1lYO344uxLRjVNimOYEeN9zC5pp4JifP
Tnp0m45e9DF3ly4qGqJi5HBHwWoNwPNlTimqfMPyOC0Oy67mURDH8tmt0xOhGRkLYIqQJwq9EV5B
C2OKrUCMJ4BZpAY3tDWZZNh+ybbyGI/K5vcOO/txwnyFZUjQBhYc2fGM3hzpbF8tLNdNAn/XUvOD
/7YTJvcmHzDTOqw7014FGo6FBar8Ho837fghYbz4peFHw1g0oPXO/bSDh0txSFrM+ARuHKplb6bA
vXXI8ptRGDh+hdegAs+2CkVDyCrs+zTnT1JMOYmWMIDaJrkAHJFQ+lYaMDRggnUDlnCA3sS9sJwI
TAYE46ROhLRJOF/4fdEb1SSnYI+xlgeB11hi2AQQZhS4Omv3W47hOk1wjep6IyAE/2jupjLJ11PY
n2czdkyJ1J2YKxqTqq24nfL4bIvOMhoDlQJpYMFqx3TvCBseH+Bu758fo6+ugq4mHmBW5dwEUDk/
RJUdjw7gzT3pUtCqKeF60SlAV49a359ShDmtc5p5GCsk/Yyj4/K7eWisHp9O2eeQA1j0+kWlSylV
/zTrh+3f9DMzr+2oFmH1pdGy0l/eAhKfrsjuo3zziMqX0nPVIROhGXbHwj52ouY6JyHNa/pcIfHq
v2gmRYMeOJrjoiB7XVjSmb9V3lE0Y/0UqNlEH8cBXLgacFySH802KlvqGmYxgnHBEDZ5IfE4wugt
DzaZN6uXxY6ulNpDhy1D5+5dmECU4NFphuMnH01f/MS48QvUbKknFs7xKPUS9NH9ns6bAQDr55Zs
KL14kQ2W3Ng5lWvuAwXvZPCoAIh+ne9HfK3u8blbM9//jroDhbyr4N/GZDCd/pH31gREZYOXDsR6
zJbpu9FHDVsBUgMAEnZScSdkJqnblvBW2lymNk/YkIID+BdJIXmd8thFfoJ8yy93AAjYlnH/AmVG
iexC0mza4xElebHRMRRA+R6fHO541RJnfth5unNSE2E0If8PJsFjeaZ7/z/Hra3DHH9ygrbQFUbk
J0LwCK/+eoHIb0jXKDwv3VzpT6+fwldTGhrX2bnfl2kAal/BJfLsCgH2GSRUslu+bUIrYQ524sh7
2sC2ErQMDTobBlygf6FgotmLOPgDeGEcS8X/NmLXuiCEEqbNRWKaONQ5Ezk464kGJ0N9rQHQVG21
efjVkEyo8oNcYtAg3ke/cSsRgUTyof2Pt27GYIB/Tgx+qQT3i4JUd61FYi0Y67WSsQv8XIv7pwwA
RFBzp6YWsUsSw/rz3+O9aYFzlJy+CCJHtdhqgNE3+lSpcSIpjcyxIlkpi91G5Q2+/zLKSuRsbqpG
4KZv0pRWJ8SiLy2LRSfyFcHD5UovbCUledjWy8PkAlpcL/ewbXVmfvIeRtfZ2nOWp7Ss5N0bRjBv
iLbW8IWutW3pvISlvYWAizpCahbdUBjWoDPlQINfRjoWv4NGjUyF4Ju5nHYLVZzcs54qkKJU69Ap
5hNBZ3RLeyMtFJ600dZq7RYi11y+R0mIEvjHjE55b3Ww9oxuMzzGYDH+mvxprYw7Zl4gnEUvxUNE
OC5WolDyYAe5R40VelYlcAe7S24STlk02dPVYmuVvRZkWjfdPLUk30TAJC88g8oEkiIy/ormUBpf
cFpUF77r3hSPokt1BJgeN8HWTpl12FT0CGZNMyv8HzKQRwnVlvrqlELPYAQY/733oQSPOrlfXZu6
MaXxeQiq4iAXJ9O/7o+dVeFMxi008JeTg4IfmWQKdd3FQSaNQp0h1DuwA79pK76TzIh5n6wt61wr
2EEQX0Knsaf1ZAwD0+Y6kMdCil/wMDJ67JO3FOI7epxkLakh2wOMawSD9+hL62/siXYq4e9v0Z+3
ad0yxP6T9tyFPtPCZWcZFmC3b7KhowcM+Z31d29IfMCT1KOddeqzFB2D8NGJJhbW5j2jLi1zvxsH
ErRvC+n2cK8DT1f5G+MuLuaK2F6K7x5ZGqD5IiZ3f6tdtZhPiNhrIuHyXq6R7vJ+xm5lAsTJQk46
e0laxfxNtbgf4ELmXimmLz7AR9Sb7LETQlb8ME3Mt2DWU0Tx8709KI7dbl8KjTaUDSYIqLHSdxzR
ch4e5yRy1fA0n9Vf8kmHrZyzEQTwCk2XTH7GCLSIacvYOpqOowur3dNRu77uUjrPd/1DMEsAbnyr
Yk3YM2UryI4z8fx7vki+le0tp8Zwe23X9lvsHgw/44+jvw8Gs9mfiRP+GODzQcVOtfqjXuR2CgYG
SBouzUAQmcAQbbzSbhiraL4Vqdqd6FumLb0fBdTqbfBT+Nn+v6Pe7fbOvrEeFb9O0X0vgaBER7s4
PwbqA+6+YXFiKDs+1aMMI1nHxa/r2G0DeL1XxzT2qBjtm7pTj0OXESI3zdWsBtoXhm0hiPPotXkg
QFprlFU/wW9Cq84TUnOMYppK2z4jK//6ivi4sLvyS/APfrzzHsAmOnrAK/8DLWaMiuxMWWlWtbWX
/3eYHGl+x7qQ34Cr16PO6Myw/BFFYCR8IV5Pn57O1ZtY6Ho7cy+L+057hFrTiYgDY370q22ui9fE
6dI1zKZP3J8udwUWTpNAT5Ep+zP+tKJsl6m15jHqujoKKah0NTwX5gcoBW7B0pG0nZP/l/UlBdr1
aB01CAn6rNVnHVOkfX8wrG3lHk46KCRgORfVrxYrusCDFF4k/FU1GSqe+L6rda8206UXNn6j3m9h
2WwPwgZMv2YHPsCFJZesmAtk4TyWsnFDsR9MsyMOsxlSxNEqrQzPV9UreJiegMMzhF9eMlDTTMJU
tah5BNGkXBgqZCAq+yExhjJbinvJj54mPCBWCWMChGIllopsggb8wV67oEjszySvsrQSY406mzf+
d7yl9smQ1k7MvM+mNAa3crwlubLoyoOzysas1fsdr+1IqRe8E6AuvjRimsoLSQrWhujy2vJdxRb3
MM3wonrwjOjaf6xN+Tz8BLHIlroL/c4WoGvK1rLV0CrC9Ixg4PoHwPLzA3N96U+x/PgR0djUgnhi
+sK0tyfDknELYtC31Gjlfip5dEJtZEn3GYELQfnKIFiqW3khOxSMcYeabo2r1hr+sgYEVySLt7oE
AWU/BkSkGd/q4zsvsDuj/oXR4dIYG9oHnsw0UE2ksqNXIWOaZ6KZvh/7m9TmVc0dmWSRoS8CsKQy
zDi3Aa5DtQx0itfjOSKA5uBEqHlT7pICTLiR6fVHoHbn5PQyzhx1eHqjSz6IQu/Cb2cDS3KprYBw
5JsZZ85hT4Kc3CGfR6eP2ve6Fe2KvH9Sc/HBa4UAyn9o0eclBKPDrBFQ9ZKDd4XxtkUxn3qCuhau
dKsUJc52Wv+peJ9C8WXQC3ya3JBRi0xMXypDXl8rXlMVhNZQbiZbulR7WXu9IfN1+JyTnhWLH1gx
PeoEqD2n0pBGivRZ1rA162wMdXq5r2Y3pt7T7yrbY8HX2zXmSfW86S1opwMXxm2wSd2LQSEQmxIi
o2fLDU7YWxv1UxLK6vGhrr6qv8M25cWUW7Pot81O0K9C6ek2WTZSxbXyOKsVxZ88y4mmhZ0k7fCX
mAoNItiOcAa2T9193+WJTbWB2U8FTCMl68eNzQmw1rlyMKJpBMA1zZg2/gxcX693NX3zFJBuMUqI
NIs3KyJcrD/GR7MB8Vr/Pk+3b72wX8EGIMKqCchOyBR830JW+eR7ZQk8UuJNyuBW3ETO6TQf3Kp/
dtgLxu1qJcVOtAbrcNz44P7QzF2aMENeQrFYNxtMhy/hdXdcZQ7mTw0C0d/eQHuzNfoQUSijX/ZQ
R8PiWErYGF+TZn/EFA3+3YFoY0Jx+uLSBhNJhESnVC+zY4U8u+cO8iRxPHVfNXaIr38aiwih5ecB
k9/FTGBtV9zUYuI/MWUCQ0VK4RjbeFXCOgNKg0K1mpMgap1mqt3R3P2amecrSEikHYG7Kmrmz6mk
hKlTf8oULULC16+Q9/rK/GWLeAV2JxyLcLRba4FqAvKw5iax6qtpFzznS4NPE2jkQoScF5HvZHMQ
1/gJvCsNT6vNNPr0vwcwTlWfcXcyvxe4P4K75ZFVINJklZ06P6iveyyKrtxBm7K4+w95prPWwR//
09J/ZJTQslJy2ob/Gxm6MZ8qHhPLwB30UwjsCzOKE/p4MaxdAWq5gWOjPu1e+d7U2XUXOVErgPi9
Iww9MdN3fmds9Jr9SZUtSAvxqd12kSVSyNda0lQKYmCNgrNvn79KwBnO2Uyres2Sfy81cGRO97tg
FbTNxwgggaU7ZrMMD6r5Nr59x/YFT/j5F016eQ4/L9WO5TRgsNIPN99F2iBTOi54CRdih3xBIzrZ
flLBm/G28462Ej0fqPSW8Xy1WHIXl8D/dQpqwc9SDaU8fuTJayqcj53b1zMOtbGrICyPz5wWXZFg
ydW04jC3J5f6Z54TqKGzx8oXoGGO334T7RB/HPIxlYgYusCtaf+6fKzw/sj5FnSxau4X16zwRm0C
UZCxf5OBwva4fVnYn0xOF9O0ETOzq8CiaKZvmW1q96EJY+tjFUHOD/78nKJt0FA26SadhWJPayNg
jCND1iOOBEfYqaHj1HbKZcx0hT1L54apOGGRziP9MD6/NKhjTX6Y1LYExAyxsCaQX4ZE9B0DfIUB
msTllyCLlfhDC2gm5qFpOk3AY9kMquqQpJT5eGjgxu/0nIA1gZLHWA2mVoLBcjDPM+FGnB/jjCBg
ECmqy2UwmoG4c0X/3nwN2xQw0QuZLld2h6Ias9MPLreusFlwlmOQ0Am9AvOSv7L/h/EVEHKBdTuE
ArZFyt1hgVXuCFippcPSV4fVwVd2STP4iEBuIBNnEcUCHA/DwUtNitR52BCsn0fYIdEZTK055LY/
wjM2+KMjgagMalXsfOjj1E7SlyV5sPlFTAnXbSN3dZ7Z0X/wYhmppxH2p302uxXoHw2OILmD1yNQ
IL2PuZzilASliLxCSXSSpAZmOEyTDSL0PngORdimMWaz09wTQ5dnQ09ZShAsWlputQm67fOhTZl1
S3U6UU60X4+nfOEwXX1gdVWZqhJvFWF4K8x1B6n6QiytJb9WnJyLy0SnvBYp6kSr3ugklsjpHLB9
qcxpv2zaCHQsAd5ONo/owtN96kt8gghRnKFfwD1u5kl+W1Pg50ZnwztSaf3+FTxVe5P4S5D0WXNQ
1WdGVIU6cH5hBPWYUN5qgzdxMrdeFMEeCv1lFCONEcQCBaiuZP3R1qpDLQ+E6UOLta8ElfAmMOvI
ZRqPCczxkRyds1QJaPZ8Iwy1RzfaMB43mEGOXiZEhkbUbLdjkn0u61LsVYVltBRrMeycFmW5dn65
INl93uM8IC2YuBWeLeSe5TBCb4R/FYe39OLO4HlkihZM4i33rKBM0sl73//D5RJNm0cI667YrGxW
4XvP3ZNXF/wO2osZamsmSE2aCKvHpZZp+uHjOMsGW6UozTKNXreyhdnOm+EkNXc/TIQLEFzVyrvl
221fnShmiHSF3UYeyFGOGHmc0/jqSVpJvpRZyrVA35+TpezBv6a1tyGkCeEcqSPha5zWhQmQSqKk
k76DII2qthl0QhjTpuQVba911hnAizc4UGoY3pORATrrrVWQBU/JTg0gm3QeqJjwTjbd0oHfEmLg
WUSFTHCsyFtNhOayUPImTMrmvnzbFHCjNtWAmSkH5BhWEU7GdmA/NsJllR6KMFvUFcCTJtL0jQvP
ZRggN7Zx6PqH7ZlvQiw2wH9Ob5gnVjoa+visNWvoDs6H2TDzvCBF2ZmewhGBsB07Q5lH9uCs9nWQ
pMUoTG47wPCCsJr+lTMJy0CwmzJQ8nT1WyyESgeMvUe0mXyCA5Xv6bzAP4lLDqEaHxvlmwcZ7NTB
VmF4oXvq3hDzbOLHX6OEMzVh+OMXHD1WBCfaL0aIwDbDY14jhfphU+7LfGQT2O9r/spUroVzfnyk
cT9IBKS+wZiJTSujyBIz1lj3N6LJfFgKV2rboxopq1nja2ONawmr1SncQ3O75u5aD5xvulgirhPz
q8P4mjuILtEk3c6gP147QGgPAkud17b+Y19u2moePq5S3gq2chlXJkj5yRmSaxCSwYPG/O6kM/sK
hAKeN5J4K88HCQwmQ/9VtugILzdKeRNQ3iGm3hVGzrGAar3XHHhjaR6XRwvBIqhcukYSmwuOOyko
5oQ1e678M07vmOqRQrJjqzFEV7te/Okn+cHAtsxI5y8J7RklCXyegJ4cULY8IzODqDpKvnVwkoS8
vGAoqdeaLeDKT6vIG8e9xObuUa5kVPxPgd/yU3t/Tol4hwxZYQlfpA2oR5ReQPkJhXzNztBhHCbD
1VMt8l6zo89MuTYO4weq8IUi2px6pXuQew8i3LChj8VvsHeUim6yo/ufIstdXD5FL/ZD1vg91HXM
QrOmUk5DzguVrATG9DMicCjNUZ6fgsWBdVaZeWS3YEFN2v932gyzki1ciFCNfaS4aHBUMp08UhAF
XYeefq9EBKxXaq/+L0tPBXu6Pj+4ej74PGsrwIWO1C948tqIcA1S+Mh0I8gd+JB8SB2tZPQXrkM0
w7bGdvLM4lATLaAAvOkKuB7To8klokD/vihi71rGzw7oI9d2JAiUyuT1gwcVSEsRvkjo5oSOt/g8
o1U3CsqktuflauY/lSOl4YYzDqFm9icU+9R3h4lIr7XDaozMndIF9ubft1au7L8B1MWoaG7UGs9h
6x4xohkxXmALo201AIqpDUH+NjvBzNic6RBekNCNXxucuptA15OUdhXZDMxqUnh9nRFQqO249Rwb
sf/GDrNEAuC3LFuQmLHHtP5PgbvERidtxS4Pa1bGGUGiyD9u8vnnBMpFLbGW/vKzcFeRzblE9SN7
Gx+Xi6ncYnHDZ/W3WDXDDu+gbcNrK+qLlRH3zAazMzHdvmFeQD3VxioVBECu76CzaYb7pF6+MVXu
bbx+V+1savrbB5a52EAJzWs8jcCrYCvIXmaZ8WjS1wO1Nip4VB+gm5Pjq63ZEqw/7f2zJVPM8kgV
l4gjuO/2jAzyzwyAN37PQH1cMAH2j4Ac0tQVEzU0GxzDPhdtfKkFbauy9aI+5W4QLFjpUBj8CF0e
IX//dmwu5Mdhsd0QGpuOA4m910LQ6XKBmgORYqyFPtXAkWXXpdWr497KHRumNKUBBtaWcXGE34ls
gdD0lisDhIm679SMgtjs2/LYg2Zb6ayt+Dxl8pQP4+YO5wGs8j4ay59HjxpVlwzyRK+NiCwjjxPv
eemotxLv+wCw18TP18aB3QaZDr1+1vy5Db6hXpkz1wOAqu1XhHe+QkWXAK/GlLRDJsKZdBKkI22R
5aGHNT8tVVnTK1wOULK8ViTpPowmhFKHJe8KBOtrGBcUDNLEYCzFFAaBOvT+64VukCQgMld37a/c
YZdEm67ncqOu+3ra9tTvT9ZfmZHAf3wn5SqgAu9451lx3XMnEX9lVN8DQfzWkQukY2UYlAyBL5IC
TyFZO7Mh0mvjlzPN+WF9xZ8x6ZG6MF9BguZeLZMwidgNYRzch1IA3f5i+2BvMnReQo5Po7iUv5Ry
V+d+97wz0Fs+r6gxft5Vune4jPZ2qUfEaFod1YG1bUy/o6jYm0eq4grIWLj32s3+9PKbmoAjxI4Y
PMOqWQq3pG4bL90rnua43ZfsCyrkdEFMhW4PNt2Q4Vicv6qda6oRtjyTxNS/L8L8uFtT/XBXmN/F
YjX7M+GLFP+3F5ta3ZG6BqxJiqYD32suvYXcrakYpbd5d/x5scpb5JtS0QcMuQ+r6bLg1jtFO6Sr
VoTwzNHFIPWTS0tjVpqBUlbSnA8cTWddh2pCM7tKLR71bCVMlwYcojANhvlJVuRG7DuLVP3U/NJt
p400VI8bKjsWDswmWvlYw+G+glJ0wzwoPL1qs4+6ZumGrRCjPMZpIAnHEZZLwiIGJAXbLu5gMTGz
k1H999m1kjU/pNpdQbjlWGviSqw4KRr8/hZS8aw9GRGU34ggvKf2Z/vQOnSu9fZRnz5LNUc86m1E
ceqg3Fy2S/5Ad8G8XNoMBHw2i527qvJPfQVjLH0yI1yq9fPR06UcmdkTL69FoJTT6d6lokwVOrYC
hPkbnGzglOr+SG3C7V3isc+fdkwGidZBgMgDUSTfMmmmBBUy2TVRfJHHTT3TTZ2bD6FIZRUtJt9I
D/atqwtgLiRB0ddrv8GCy9rYu7k2hEIRqmsnGlF0DljEu6C0L2Qpxg+xUR/0saIBiOw4i+CdeChW
ht27pQsUhfNmwQjTlABaA1c4JmVVMaVEqbpes17LdQEt6Q3/DhCyGPetf06MupegbRRerBpqQIvR
gMjfXN94Pbl883pAE0RU5aU4dUULDPS9og3tNHrzOIOI7rHc3isUexP+thDRWcSl1ix33KwsIa5+
gVLxmTsWlBg3QpSOBGWbd2ypxLIWrDpLt0sOGVrIEajXKFYIukRmdgcg1DmcfMtHP/jVBINXt2nX
kikIHpUuBGZGW3vJ8syrkKDnXxQN3FffD+7fdm0v3wv/dd1aAcTLlR+KpI4hDIuC1ZoxJnCPwOK5
Qn6qnCgAKX3ujKPKn6gQMuCuDqz+sriR0s6M3mT+FgOiO6aYoqTA9ZZvbqOu+icKyCfmGHTAtI9v
nFw/JPiTvwrNp1iNoNas8qIaVEOkNX1cr2nlghoKapeceU1tso1Bla/sxkUm/wqmO85ljC/dbTei
z1OrYh79WmmVIBbKQLmON8rXOFmew5dK++l7WwGL+IFH6lyxzAcWL6SUdjHh/ht5AyGq2jmCgjR5
JccbAPHM2lzrABAug3dxCNc+UliBAgQzl58rwqlW9ldN/t1cfSB/1lYHUh5APG5A5UebDrkYuFmF
pgB98OT3UKH53s+EnJgDG/WIAf2B9q37tTSeXvRWb923Ie0+0veLobSfGhE6my8m92u/MBpkdHao
iBDJ+fDSOI6810lSJngkEDhTAE4kdcUHQZbMZ4O8Ay82rpHADOtHSoP3jgRZlpOtnXdlonomaV8T
iR8N++qOYb+hSq9i4s5VofR3/OBAYR6POxDgI2qyQy9k31Ca00TzBjrAd7VCus/MOQl9dtVk9Lc6
Jk3qD1W8j2HinAVoW9jnq6IUiNf5YclW4g8hcW7yF9Xqcs4s8wOBv6o7TZTsAjKz5ntEBzxnTADC
gD/nt2L0rPOrYyuaPr+fIZmFNn9xYww1DXDlo2wzKwRiCP2skFDjPIYuzttURehQKnuwpc77bB6J
uRtCNJJHCbQGBJDJeIne49mApMKQ8A36mM2VpF8bVuWo3IqRX7DQEuQl/StPYEYyccdIvlhYGtvG
aQOvbbdy5BRfTSBU7OJ8oWp55j0vGo+hpII/3KPzPAupMMLx3g51lApChMKhnGPFUaWbjJqt8yBn
YfutDSHi6OuL/qYUCSeZ3MRHn8DW6B1ldydEFnQnl+tHhhwJgA1fYWrZL2VM+b2fPQZ1TjyeQ7SI
Tbj6RlBaAkO3K0R5xZtBfTlbu3tF1ydCjvpudyPW16+qVRhSzNzKFWHwtMpZXtlm3GYHszZN+lJW
FOAaneWVcLKBDTpJ9eUZJJ1YV6uNcc0x7Nw19Auf0m+DEk+2Ghdk2nG3M4UaUbmGMXtUfUYEu7XN
EONWNUnMqvAFvsMKqkli1VTwOaflTe00+0K3iGUCUOKJn5vp+U9+vgTCosW36N8ZB5RK22Vv79fP
G9ZELOUF+G/0WxFjnEFQy5j7/nEha3Tp03irv3oUH0Brj8xJGdzN74DXX/+zztkwTryszhppIwAy
BCa6gPNPGUMsH7Tfhx9mDzxk/JH8UMFIPsgkupVIlD6KW4/DRBWoQAFIONC7F3Kvkn9PmQ6i6mJt
JFx26rHiJW1WlmiJeTKRLIllnI0bDDq5+mWKYJsmhS4odAC0NKuD2qB9mvEE3csnDjtFcLdMt423
k/SQTxz7jhK4yZmCOMxmpSAGOjFgreuUDUKU1iLvrsS1gLs1+mlP0OezSdPZpW6g9zgcT5pdKUo6
0qmxkFwEZILjNaZ26PWgFKxnkGZuL2uyPM3sa1oS0kQ/rsO99s5+KSAN0BIjImw7aGgfXJrgiNw7
wsFrmgm4GdYHNudHwbPEInCxFaB8Zr4OZgXey9dzKg+nbW5Ht3FvIB/nmKDyjdaW+zhAX/dwpCWk
dI8imMiJY90yQcME02jD/nDHad9/JC5wPP/oIW4NGHB2P8VFwoZslYLFdD6lSmfYxLvE51s7qjsK
cp4E5GcurcERpe6gu1avcgaZsR6UXBau90GbhMT+FQG5EL3xZsGQmktNQEfzPIfiAQg2gmhXpvsy
9gNGpnY3vX+m/GRcfefOoJh5SaBRoW/mVNzVkh8vlKwwtrDGjk0yAxjLMetWcZrc0fvFG5fv/oFe
SCyEONqH7n7TEdzjtePacfV9I9zPAigv5nbSXTY+RHSxiTt6kpIDXEdNaHyCsI0outQuT+0BzlF4
ZXkIEgsreigw5jTVpy+OMTx9JOiJLcVKKxRGB8WzkXzP66qIYbFj2yaX/cJ1hZHmP1ByLL+uCmNe
x7CrcqZlrLvzYAf7d1azUL3yd68WFKEG04n7Rh2csCJWzpDjKIMqJrBx5SEVtYifqKOgccihbWt1
age72W627AYDqS3Bd0j9OMnU3k4S1BOUw4fZq3/s3hEHjezNEMeLUd9uBW+kIB8rxeKDlNXKxTbw
PsbkUIy3oFqVwKKKok+5xhvZer1UkNXxpaMbQrS8d/E/uerqWfWWUdLkAEEw7UOE8wYs8JcEnZs9
Wiht4xtOuNHSGi+d2HANwXKI7xKlSx+EYuvOFSNm48Iu5XdQkfl88axTuGKylhLO3SaNjTrQPBkz
9RYc/PlYJHOiZ0i392j662bBqlC7xPEy60+hz7tQ7xNH8kYs6p55DSggMhoWZemVw3tHuBT47C8P
+fYD1jE9IgdHmON8XDVMCIWDFWNQdAN8ALEIJvzGT4aV6BhOzKB4cvsaX92SWldd0nI4/x49f+A1
mAIN6izJjTeiHEdIpELPpizJTUxPPGXoCabN+HA6peLStxZxV9sR+2etnJW4od+8EvniX3Uc6EG6
jdRHMoad8q2ZthYPHlLnDsA1iCTneLTwVIkzXizlUlhY9jOxbbO1Tfftwm7yoJ0KUEwmfHHURR+l
ws1Q1mZ0C7pZoMlnfxCIqb/458edG/GOMxDvbMrDRXx04Qvqgr63cDRTE7yzhVQVRGDK4zg9XUVj
wptJIn3yIkR+A7nlW/F4SWSYekv8fjNEaAwp+itUEAeb6ryub+RpxyiZmtHh/49BREq+PDuWj8Qd
u61aNUYOo9xAEKY/RVHsgJ2v23qii58cQW2bVU+PXWalcxpOKAXe8uqCBDfzTGxkAyPNx7YM3g6Y
VhXjGeofsj6Mek1sGeryg/EEh2FXx78Q4InRaCd1+HTXmZOwE9GKaHBKN/cIXOCRQGyRwPB7/M8S
idNUCqs4mcYagESyq6gr2/8wXZyorkHqkIjEgOzkPpBRq3gIDnRQufF5nhtMeXXXE++mr07AqrVU
uqDCR4eNCfFPjFTpN2eok23rbHARnmry0RST6ZwGijOMMPq93wNdxrPv+Ah8sAVX8Tfrg0Qg0sX1
UyjqWQkl9R5t+L0L03bUByz8MebIE5+t6MylMNGH/rSIB4Z77mpPxZT34QfrQwMxUezB964OToC8
PqWEoIBVtwokglhnIpu+9RHktNh+LairlcSXZ7c7S5C+b9tU/CJoT0FdsSVuoYBdfgasHBqwZcDX
RZa40/DPSz/bSAx2DrMOp0WTyqhZW7V8QoO3ehnUaNFppnv6n+s0Y1DfkP8ysGCMod5T5J5Ut5Of
8QICzv4WGFNMpLMLs+ew51BnDwEE38Gg7jaYXC5hZFud5ptLEdrzg8HAlNQ2fRezITtSgblevlBf
1DrFcp+2LqkC42IEZ+mVYV3JuEAUIG8D5C7GmAnClf77CF7N6o5Gring9/yEfvVnJtqMbWJmKfIL
37qwPJHCQI3Sna6Skre5LdHrW1R1oOIAxwmaaakbEWnXnQT46E07pNC15bYsk33WHlPSm9kD/UBT
L8JhL/z2/bfOybQG15pPuAhT4ufp3NgDTZ3N/M0MPec/s8Fim+GzWpHT0vHlGctu1h0TCreqFezc
3ppt2aELYoP/hKiH0O7Hra4OIO+RZctADV8D3hK3mt7LWyGfIo6Uem1rH7Bb9S19RfLO/x1IjFbX
NVnV/bn2QnKyK2wqFD+Yzi8ChajM9URCplAoVYET6lDVskD4+kFP9+UbniUZiI30wxSnqFyJ6N4s
0+O2ZvSX2jX2nNgm8mj+e0eS64l2nfYZiMEVdMCAuhXz7fepEtTVZ5Xbab4zy3hKon/gLBJj2cVE
LJSQ5/9/fArkaViAoXLjlqAWDcpwexDLjCw0fUW9aT7L75cHzU/fith/atTywFVhH6UDRlkrlhfm
gWpwLBpYJ2+MWnmtCzxEEcLwzuRWzxd6U7wN6FJ+dGk5/nNzWrZX6qsqX12Vrne0qsMXlaz7VgMg
NjjPBYeo/B8+AoE90uS5+1M91pkacr/EZ0egE6/w0J0ufh+8cSaBWEv6CQoBF56ziA8FnbcEzrBJ
JBeGzvYhxAA6s5eyDOVuscrBMMOCoJF68MDvbwYMFnsELrZzH1NlzipYVzaEpSV815HhLaV6HaYJ
pkiKvGmD6K6xI1+9UzT7hpf/jj/S6RlwJKz5V1Ta0e7Cx4fjJO0ju7xqvDwQunojuOd6Iu5n66Mx
ct2T40TmYDBUsJCkIeKUJwiH5lNhoCF0bvutewJWmjWTuwqabZGKD7laUzq+8j/wAnkbrE8umtU9
w5aP9iB/VUap2/htZo1RBF3ttcGpZbAUDQuSNzw+IJQfEj+ajAh+kbtZMtAS9Dgmc2jJDcCXhz0u
jz71My4z2lK8mpNBrdov4QO7C+Zxx1ibqWwPtpysKrwCJJb4yopUJD7wFNatZRezJQ/ZuhgIUngI
iknL/UWQuFC/OK5Q3FIGDqShZJf54qr7o9FzHCrG1y7pISQndlDcxo6/87SJdV5tHdsdrMqh5LaM
MNtljWamViOXdpzLndyX7MZuJ3DeltSVr7CiguqgyjA8M3DHD8iV+XUsNrGB/CRJpm1892QejjgX
mm13hFC04g6SzOSj5J2IwqxkKJLG4hb15BBc6Ca7ixV42B6AH7lcehGoeEUIL+VoI32cNomvAs9+
Ue6VRsnMXatnK9+qkWHOKgNRNUit+3jF2Mq+644Zl9r50zgFwDmHqqz4GbhG1uAnERF8DKRy7rjd
dfnR4314TNrlbIGB6dXYhqTodN+HZLIIJALBehX89qpn3EJsMtqIWPbxvzRIMOxuqKOf3afOvBbM
qecClOC0eMjW8ymfw3WcQg54ve+7U7cQli4NUCpXuo2Kvm+uAES7T1xPvo1eZ5ZaxKq8Em7u2bXH
tgf78c1LcbBAiUn5/6GI7tKXjMCS452bKuWo/hbcaWBpcxfduJvVVRDWnjygFreZhAbwrPsDIWt/
XQoQEjEvj8C0FdqJhTr0qOwLQHrTfJ9MEhW3pLMPASkBerFkyHaY0TFpO4VtyI04pftQ1P9PoA0p
iBkH76Zi3Nfj9ZgpMT2C2RzEnwVaVJBgxpRO1MoVWeNKBtTch0r96z5n7ptQslyGOBUdqO2NSSsj
iS/z7QCOmbQVotLMot1fT6bSjE+ZjFbaBIoKAy5loOdWeAck83XKkPWXrOipVB41SFfOvPKpoDXR
Y+2YogbDtGra3td7hQZvW73lfv7MZGBRLtMkyYb1aBXb9CQh7VUAiisDAJh/nw/NAdEz0t/zUxe+
3ag3msIjYxTqJtzEa/fSMNtMvP//9sMWZJNx28a0nwEaBl2zwpIFuJFEwA8Nr1uHexheNXipS2Mo
8e2eUCu3xQcGwwnlTV4zk75pqs1C3zo2FAbsjETMJZuz7bS49pDp+EioOFyVW0+LIKZAzQvZE78X
PRQ5jvVK0/wLTkBaN4VlyxzvDU7MlFybQCwUzY8cS2A8UWvQDc+tEdtbc0Zgq0ZDBrfCfq+n2b82
2We8iHqs0oD6DebXh8PrPVSPcdYLJ633RMKp00YI3rSYu6Lb91Neu7+Fcu/0rd+uC4rUnK6BPJga
m2oeZnAxBR6kZeRQcoRMsCjjMfASfRF0lUHai4dh1d32PiPLxG6w4iMYMwbi68pRItX/X+dRkTvo
UZBQ4Fu3Q7NDECqmDVieG9osN/efRpEoSfFLWcD5ElRppiy5buscw1dWFxR1V1/okX5rb3mfX4Ai
JJ7DJp0n7YggAy6ljfVBHmyxFZi/mBIjFjWHtOGvl0v6zK40Auq3oma2v3I463eRuBG6oU0W82Uy
+ZW4CuaGG+NwGH7BzTGNUuyug86mRyi3Di6Dp3Zk3SzK//DOdDSMtAOxWMBpE4M6KXDVWvoJRkEB
SaM2P5p6f1viwmaWb28Eh+PxOnSkIRk1WHh0Ht+GD6TkteGl2QVprlreh5QeAfYi5R2xsRwKdEJo
SnVwCfl3fH8DrlrP8sfgW/QR4OCbWsnUhtmuCNGE/n/L9DgE35bFmTRst3Vywbub0oMEmk+B3qka
Nxi15DALeuSKUCGMBShhjqYQmLibxhQDpwiPs5vvBWQcurLZaY0FBYY3ph7H8M9x1vC4ICrv6fLI
WIQgosL+MjSOWJfj414eecHwcmnq8VQxRMEMm24x4enajCAzT8LR8/3OqgqBq1XFBJe4jeEgWaqi
MSE4YfSeBBdbUSRbdfPbeqY2jSNBtq8X8rAjJ+AMw6+EHYnvCh8aomBVtOPvzg/WMmmHWmgw15gT
5NqM8966qv9MMX7LoqT/urQi3Kc+s1CWb3sWaHVMyVTpjLZdBnD1QPrB+hZyjkplx/rXNPrI7ok4
IOJlFDmWgPpA4+vRpgRnfcy/PHgNBAHWHeCHRnb+p5ng2h6kr8kyt+931TBYVjdL5ENy7bdMnZ1W
5MGKGyLlZ0iVZ1T+cvVHoKccli77ykID76w9REoTs7ePp/TKNmlOs/grAY8Kxqo/UelLZMCHYXFP
EVoPHdwSftGzS57EeTehWTtarenR69ix5WiEgUXOt5wxbyo8E5U66PO23t0Xc2RQ9QC8aPXnQ+zn
gMeZxMYn8Bw82XeEdd7aAfdyfxwp9CLGk3N840jD7SXckWgXIfHdhHiwdsy5H1oiZ/z/VQElTDSH
JPQW6gfG6kudigskgMQuASp9HmzCrNO+CvGNbPIhfkM4sw3rRATP0vK+ofZsJGMj7NzcwWblAwt0
F70bsXd5clP/t5MUna6PN4kHZrCl8l0769+zI+q7FtVrwvHD2iQ46L+j2gGRiRckD+a9cAgQIlo3
VaQHurFXWwHfIIz+dqADtW1hvUyQ1pXhIIOOnm99pNTzpMIuJWUOu0lYCKFl9a5XY1ORjYRiyHXk
MmQbyJwdNzUs9QFc5+jNEeIJepX3MrosXIQFyUvzkVzGjxYa6/If+wP3gpuHWGB8QIqbn+joi5t2
oDqoayQtaJiL//z9Ornhpg9rXsT+PQ+zva+Ytysl8WytCrZwh7wOQmLpQEg6hGIoF65w/8WMxsFl
bz0KHawnRfayELBI5PNY/JiFt+9FAUJAf1iR2INQZqTjas1u/7fS2uAmbvNB8s0qnpaBU+o09qNl
975i/faI/R79RUpVHCp9yQBI9aTrncCsRopA0MZbP1zsW6KoU0GBk23YZLwVuepO/AVZ7ni0QN3z
34tDzNZjB2jvaT+TKYzreIZiczRn9mWfz1NmbeuFIZofIV9ee0UUuQUrfHM+txF1tJiR9+osL+xU
+bNThYZoyFp3kPKsefBiO17yeTxpMnjm7rhbVfuIfKreTYi4Ug5J4mUTejgkgv+C1H0ssptPQatO
kDl5KVAEbpdB5f/8tnPTABErrk57VN1iKUNDfK3qUkpZhEFQkAErlCSzfr+BNI22gfilSk54kMu+
U5g6Ew6QOeULOMyHz4zPBwtU5T1atEoCseF2bKfHXsrWRlsxp8qR0Y955v96ZWIr4c5iSBNLXdkr
bws6+N1PTbb5voNQlMvG/d92xC8Qo8xfN0EGizcnhG7/j0X53JbV7ilSwxFNMDkb31IiOSRPs48R
on49G9/uYyCW6MwMXswP0crtDh7Bp/Giw6nnkfU02yGpX994KwssdZb7aQHMme/T3JsmfyMVRUiz
+96Un6UdNVkI0j14w0Itftuid5C4jJ/XzHRo4ePOLmJC1BN8V2SjtervkbKlgvt8tAvTZBH+74Lk
IOGb2DliHrnmr9mKpN3mqbmAaKhu1rST8SN9Fx4QQvwH60SndQrjfbxizBs5tg3ihTsz25BkPDP9
wZXWhpIwYof7ZDHMLoNoIXKURdg8bezisdFFaeGEx76A+EOifwPbB/umyoLzZR1mJOcNE6l4ckKX
hWRDLs+oal1D02bMWXSx/epqHMceexuymZqaY2pqXjVgiI7FawJ7lsvl811yEzGTWbcSBrb4ZsSa
WgHAePvjIptKJcYqRB/IfmcivRsuJtz0/b5juoJ0J8n4cyVeZ0+SYsh7aT7jfynbt8FERu38qPWL
isWJkFh6k6cXtv36if7+EultHWC4g6c8zEaL40NgvoJCHwCddUkQHMHnyu09aD3JKfuyV4Eyk8xj
H+saex3YhsUe0a/aB6lid4JfFixvLa6GFhEow0AddCtiXMkcMOv0+fXe+TO4jBNJ1w1KUXYa+9Pj
rdYz6/dsIRNsQ6+/LNxLUifU2b5fgAH8bEZuPOZgX0sL1RxggHsE9d798Ls8jc5FQSZsyiL5Yc5u
EzZuZykFr6q7UGHexCPZtoorEaqt7QCJP4j67dlp8KvIhM+VSQi6dQElsVVECb2O/xzW8AUnSQim
DYqgcQ9a29IZQRI2lcqRD77U35JqiIT/0Rg02pF+4o+rsa1owtvCfpFL8/UkL96PJu1uBYTQesUt
CWeVSm1ee44QPACfm3dgtcYIvqBnO43GHDTBdygUf06p1+64pSfmvBWhHpppTKCDSVeqg3aDY9Ue
5zTGxPgHrqxyEE8ADgxVGenEhnk9FY+2pdhrPyod8moS4Q/2a/bZ5Zmb9226hTC2Ix3zs32rrrwi
jNfANpMV5zP56q5B1WiuQYu1xVaOIsLFrgmxTm1zJM/YY8BJtTWOIw4D8yBu9RPtrBVafm1kxTF1
n+hIEpsLKKlYVJvGXoJgFkOfDORfjtMEQf7lIw6LwdazO3jYX2A3bpvzmgM/58Dw1ySOAAqBRvY7
qg4/U5J67mlOc08t5XsZlfn8Dhkg+r/yFguV+JjOmaq2V3Ta8BnLr9qgvyVGI+8vfBhySrw7/vgD
jOu6BB2N8xufm1Ez+Qm34duBBfiv1H+YS5cVe4x6e3D7E09T0arK5I7UG4iTSPQr5d4g/7C4U5bl
3sRa32Wrlf+zJv94xon5bPlCcZj8OVJGzLCXBetH9/M7gfPsxFnOfW7x/9O1BTahrc7WS5iIb2Fb
ZZM8BFsQ/RPudERGLQJSbisdIheQafXgpmficf4ArxEoFoYIdiEZAyTiqgCHblSj9bzDJtZulGu2
pq7MD1LdrJ1wiSF0AKAJV7mwMRPBUlqK6gozSlbY1VAHgezQddijVZyccenSB9zCBW1L137oKUEc
7p21an5olWX1Nb+PMGb6zfnIMQO3D3jnve8ar+EOMFJoEFkWDoveqUEoEbDJaCNprDVsB7KRskVH
twL5dGgqQn3VaZ7x3ZvoPFCq86tKsch96/qq+I42psA8RZ8a5uUoKKd2Oh8jif2g8q69/k39C5kZ
t7gqRlpIRNUZZ1iodfdDOb0/orTDrjw2NWTSrZpyI5I2mgZRwtbzEzyBNEM+hCZccKQVdb4BA4E1
TfeSJfOEcyZluOtRYrD14/x0Wn25o6ufHuewZ7cUUyFs7ci3iXXtF7ZPlEdXCACaMG5N8wCMyzCN
EkyMZ3mg/lvR/1pZOJiKXsXEBIMPCx1QYK54x0fXTW2Wm++4hFkY+FJeueYsnrWSYoRK09d0Y4YC
Zfx4HZLk++8cDoco+kVMgYSTo8PPD1/HI4OOFs7T66uYUxVFZ4kJtYIy3HMf+3sV0kADRhtWPWpP
rdmkzjQ0/XYNRy6rXFufQ+DgIhg8RiOPIwA+zxMNTbNaVSCXuEp0px5BhdAIpbvmxE7Q9iLCoGK8
9KB5DPy450IIdi3zDULuLvPNkUjTUEWrRxS8QBGb+QiVglrwyb9or5iD0xV9GV32d+0RUdAsBGsK
bTk1MDM/5TrHuewrGKAwKbVo6rZg2QfBZEpVUChBtBvCMafdI0GECLgm8gKx9cEDYebHJuo9iJ0g
m8aFk1TRedl1ydDepdUgXosUfVHKAEWIUhkRPis8sp6U9/ghBgo9jZNXRLu/mHcctWIfC2KiA0eF
yrf2ErPWBOTa0nNdHymd7oFAjsWsPJaTQclpuT5KlI7ckFhoHOGK6fU3ECgZdVEl4QDU8bU0dky0
ZJP9QpFcn26uDDuLn80p1HfDsNGbIjt0J3aq+vIk1e+v8ErSjZJ3nPPd9VLUy1NoapsCtR9EjlJU
fuL4d3MJ35BepKlbDceDTd4VJd6zd7Zx2ec95WYkL/kCef41J9JnBqnLkxxxmgKTq2IWNiapB19g
Q5DugyWC500hb2s9DQlhElQN5lRewt0lhgE290AQ4Lpkpibn1plKJTf8BpcPjD+AL/DpBbA7sPP0
t1NnRHgylNlgK2X0ZMblfioxMnwOpgJnL8i6QXiAlYpvqvVmqDgSOXpTTZqMlfSmFSdwFBqvtIkk
HELzc2txxbs+S2wSw+rm+q0r5d6Xyn2x6WSLeV3JNSBolALIendTcyMNoRr1lJUG+kEhT4iOsUwf
XfivX+vbXwmAjr2EiVNM44hvoxLqYL/KeyAgzbsEq8gxdr68aLXNKIkw/FydmRtUiewEx0YJyYIN
rMZ1Z5MzA9QHq81KWulzM36iz5PlZYazzN/6c1De12xH3XNZziHcHGwmrMJjn3sZZLKR+2T/0Pqm
Dicqvmo7qMkrNiEbaEvZlNSunXS3qxzRCnCMmuPGAUjZDwabapRvtH9mFQY0xITDuOA8CAJVclBa
XAbuCrU72NUuJXdBiAzo9HMfjPjaEDvKYcXSf8/IA6GSU16bGQOTdnLoiodpYCbl1hcCgw3ECPMP
0WrqXjVviVE+G40HiXg8sOzbGlw6TYk8FA4RLlOUqI7BKczeh4vKr033iwn8pv8QJDpUJIaZGI4h
Gz/qIlRecbEyp74/YGurIPxd6YS3fPIeBh828SlF8j5yBN4fpIif1Zk0EQR8mk7wAv0ymNERxOZZ
kfksOzvYEyMPq95WYJvQkeywJ88LlmRlgc9WoF8uG/HzzLdlovlcy61+7MKglDJZp2QAruJifwKL
eUYaWgxWyGB0y1dEAk/I+3zLh4LnoTXA8t2KdK7Aoqd6BVUFj1sedfHRUO9oghVtOfPik3jJDxEc
R4IgU0RzLCadqtq3KwBrNkxQEeXiUozKChHvcbxMmyQ1Hfyob1I1SFHXcT9WWhlYB5ptMKbIhy4T
pvpwcjhIw73hNXnpq40rVghfBN7tBjCb9rbdn9biXm6cxnAvE3UI+0H5rFP0XWfUH6nAajwFG8CX
5dzpusT2gYITSHXo5cwFIvG/tANTqVyb7+0FTQAlqQJc4vAnoobRToRl9wGSZpGbPHVpSNZPk4Lm
UKAaUsWLshpWbEJKpphVR+vCybzAoyuHql4rEikOvzEwqDukZOCuA93UjQg+KYegKx/2LHu3fLCY
N7zXdPp7EEmnfe0f/G04KV5u2kYn0rnSwLMiOG59f6hlpqz+PXTTY5iv3gYa5wQCRNHyhiL6nd3N
1VwWedVtoWFxiRNQRypNRkVcwUtbyWpMOqDU7xqOdTkM8/Iz1qFm5eBgm9BYwuinqjhuPapLE9n9
XfhLJI7GuiqfjTvAGvSrH0o3/lV/gsAWhskj/1WnnK8YVfaOnLjcZJP7xVf+dLgAs+/aEssr/Bm0
wU2Yen8ZMes42ZFZl5C5KjeO/csr9U3CSPuL5wMdFsObUb2dHZGmIYS1ibJiNb1V9YsgEtRWLBOG
oXPJ4bsKVZwZZUMDJ7eYIpXOmPc9PMFYyuOtthpW+4iwtXEhWgqvz0XtsE7bi4FJzAxgKK+UpIIN
JMgCtsgDNI9fQ606ALhLVIg043p/eRPASXcQWu1+sIYcCGmD9aFyuNYAlWeqmzGerG9EmbSBDcgi
pb0cnp5HAHcbPmTV52hLsa977lhzRmi1Ce4EltNOKHPpGAJ4P8Tn+vwjN4cOzYBlvxK6AzkBlL51
Ghr8q4AFOAo9saVGh8Xaq6sonEQmZqa7DFTk+9VYZYwK1JSKgSM1U491eyt0wsCQAkEyS3+i6Rr4
5szFFlj1y2L8DZIgxVMTmUQem8KMQjiMr1k5mryv4ulkoMmvSl1ANDm60ffZHUWbn2PCcYIzJ3ik
LU9fv5WuZWywpkthA5h3iGAFPZzlljmkHOViwqde7lEBVIdg4GAQy4uVdtskp5ZvVvYapsEly5M/
4i9Ll1nh57m1QkdIrOeAGOhdFZO7NAgV+rgVgAgeyX9AB3mD7pD6XvVPk88kozYgfJEcQSL8D2CD
XPHe+sN0Sk8ZAIPmrTVqZCoKjYXk+tzWs2JV/BXToMd9Jv5pev1kwtspiGfwMFSFtItwziEe8No6
3GHJfm8JvaGnX1q1HQA2uzOx5azPlI6kky7eTlRZ0CxLZQ5iX9gefdTOmJyO0Bn8bkQBVKmhNPAH
y07hUuToP73abM8XC/5omBrmOGrEEpAOV6vGYR9clmPHFUdH+4Ffd/neLIwKzOZCGInm8BjiLKjb
DcLYEzW+7ILmpGT+K97LBXJVpCENY/bqlWt4CnDnDw3Cl8AnSJr6wW5zR49Bth151zPBKQlWQPYs
xWi3vWVIZ3/iTbFxM1BNF5vBB9vMJ0blrTHn7gFWD0g9eOeDgZfr24CQEiH1XQtJsO7rmdkXmQrc
xrWXQCdcWuHikeKET3EqIOefy72aulj9YRu6/nPIi22RnrkkXSk+hBmq2o9puyc7Ommi3UbXlDRT
slpICgssniX0ygv0DVr7SwETxfVbNa7lA0P7vueXTCiKTtYSTPPzCzhX41JAS+hfXMmD5CcmF/e9
oWtLqDBywo/DbDow2RqYDPCa+uet0nCSOlGiuDv2j41fwUd2NxufHVwBJzK+sORnz5nSr6jQUaZr
TxlQOcBlaj0q7rqQtpTtmVYh9c5qNikLnnLtaQDRUMGyBPDtllNEVfcUr0SEG1ZZT13K2yFnI9BG
vJt3yS5QWzQ2dk2VKc2Xz/uqD96TpTHvwEbjckWRqtXfhkZr2HXp2aijo5OA6yyKyKH36Ez5x33O
LE2o6sd43N/k08gKokpLu2ek/LsuwZYcypdE6NlR8KTE+hnDOytnvT+NFsJspIWml7baxnFk0hHA
fnvpGV4lfwldH1xj8oLikxbPsLkHx60JYKZvizoIz2X8JU2vIOoIL5+8utlesNfseFv4XyXbFSit
HY6kL6vVolRwOf9if2S7MjCYvEDypeFJU1pSWVZqR/+TTbBfzbH0J7/Xzd8eZT6WMlaAN9kv9ncg
QwNR4FlQ6jzByYGGGE9Fh9HL3qONS6EGryPRhMDXiFLcmPFQAq2vggwpLXA0TXbjc/Qg5cN/tJ4c
Rqsr7NcjJFAQ4I47pBuUWdiQHktoMibUStJdbNJyBOTErGFTsdwSLn+y1SAB2DU3HDN72mbGvT5x
3Bf6XCnOf2nLuY+7oP/M7DZZe7zdrMFyQxkNGxEux1JFIHNOEvIpGwzC0FTHhjx+EuFWFty1H+3V
8EVaQgn2YQVJENtRRyd9X63dT/Ixl7//ktZEAvs53X265l+OtQSUSvG8Q7mO4u6mqfNjqgHuepGz
NXpWnGATQXbi7/Y0fo+lwMkok8XAlSbPmgqCZ1tGv6V4tc3N8XhfmWEeD+HWf18moX8cv6rV2vTt
UTV6BrRGpGIrnfpiJ6b+4B4nl4ncvfPU5jNtQn0gT0R1W23qLFAQEJ8RI0mBAMEPC9oQHpaGGC5+
P6Y4ShXTiigSn9/nzQ1/CAJhu0bnbIPhBZdLL+S9nrIErSWBThmwjOuTYZrUToY+UOknTKeNOvx1
CaeBFGu+v1TcMrpG02cNHcoaoswUichxdxuAZCWrBxL98Nv/PhO1kN4AIcO0rSJAhYyKMcF7i8+h
cWL7aORB/TlwusHQNik7xw4N44N3jEvITPQCL5MXpxmiNZ87JBy5Q7wLNyYjSaAH3MZ/tyTwJrW/
62pMcG4h7mrqLRFyBQhrvCuvfkzC86tuWFuojV3jUdkmS4Ep99aYpSBaL2QcI6Sb6Fp//DJAH7+Z
VJgFhc9+U6E/kNI/ogwb+Cnj/m0hqbUCC5KrfRSmJxMYHQdLmHaym9hjMrDcPjTArrm06xd43amF
OqoxVTq/JmTOTc16+dIXk6EfDk81Ddm/clD/RhBQ1QlRBhGPrznnicpmVd0uilR5SD99H8z/wYW1
q/+zvegTJAySWhORgcu1xZaYKgO4r0+Pbbaa/IrwEBdY1NYO5n2wj2+rw94u7YFcCTClRX7kAOgL
YB9qz1glKO8IrdN0ZBjnErFPd41hqnBPTcmfYyFDuQvecRMZ0lxFGj9FllzYrI358CvOMUiAnxi+
Yb7+4dAxAf8YrzeUNxq9dilfsVF0JzOr6BcQB9Zi5A5KD0TLOKkK+sfuBjK7bdn2japvwfN35zFq
RbLms1YgTVrDIVJHViJgLxccv1G40/7qK1SOpQ3VsGEkSxy3vdhcWFJVfqaEfESAjyazbrZkzl16
tcdQWzRuZEFARTDh7v3y6wX/I7V2CYVxW5ilLN/LYfXsCXeWOV3tzqhgv3NMuLW9KyTKQdKoc6AB
fpuMZEsZ/LUAsa6SG8Vm7BCf4bivQo3wh3P0CeYvDgPqblDk5f+Yt5xznMNb/j6t3NmBr7tXO0FI
S/Hq0oE6V5cnNUmHoa2P5zwrOW8+Hl+KFN+kRt+uC6wdHx+JMoGA0r2L6YNc3l/QQsJaVvb6fR4b
q1KoVDmSZXaO04dEAdPH7FIgT6dGggKzZp+zprDQt7QyM0EM/jjbXUHqne3Cb8bQT+0Wm18JUnqw
OBvF9a7/LVRqX+c7lt1UhJ5H6IaqAJhKB8tG6xx0IisuS9sPr/FZOqg6iXDYVP1CutJun/hppCBq
LpWwFgWdsDmRVhk2m/zfQVJSNPBSF2XS1I+6O8i1UZm+s0vPJaCbXEtYcpKGDqyVO2sV2wuTg00i
yQBLQtNtqv/2oy+dvGMO1LKX/z1Tbq/JVZHustMAEw6uFhsrMDU7dqhyrs+IT5oUUCHA6w7zKS7g
74QBKmVC9i8zIVU1S6L2Q/BF+ynZGSTaGpgkvwWX4KvU/96SdBZ1jK2UmwHTUJ8ApuA4STpeAkQd
yWFGYlDJ9/iIb6bwJzg9/sTTfKact7FVu6jzwYbU0WgD8WAaXv+HFJSQAV9jQArG9QyunPU8K3K6
esZsEPOJt5f/c7sjbd5OqSV8gbahD6Q21mBDpe5INP61ci+VzaVkgisGjH1R0FQVkHTbaFspbyVP
90dx8idFa7of5xH3ibBV/tSO8PyyBBtVBqrCgv0BAaPlBebYD8DayKtdaN/j9pOqw8F7l2SC6E5F
qb2NV9wljWPZeIEHGY6sMqshmXG2CLsQEn22Ncy53W/IhAP0ry5kQnW3s1//SncEWZbhH6NmWpTs
mNPjKh9duYo7T3P5NKf5T8eYV3jSOMva9x2BXh8ICqlQe+ETjvmBjnJYSkhYllbPSJe9PevPVZIT
A/AjnBjNvgS4uBReuFpCpC3mnX9ihAc7n99Ku7Ga8OJMqKysSm5ZY5TZiStqh/qFsvSUd+7ZsxCH
vAlUK5la2hi3NVWJWioJYwc4XV+Led/unqZV/m+gdEUaV+YFBzsNH6HSrZMurJ+WM2NCdbJIa459
l/iixjpZ0994dX0SbvMlS0XSF1yPf4FOLwAmzWppa08zHLaLx6hQlkzgO9Yd8RiVOich0abXqPHP
jO9Ys3LorS53bOlv1A0Or8aVTGaTMIJUisEpz2ke7kgVnErRpU0TI+o91bWo/KhC9QQpb4sfJ08v
ZGgQcSe6ZtRjL93ipGvzgjOMcGMx2n5pkOaaEiw4qZL79IPsLFaR0EwvE8/jImAhuRAkTDIjFWCo
fyaEWXOw2ThjuOUj+gQt2385TL/EtRJ3lvqanF1THVHPfu7iCQZvYtJV/Oj4vOgH9v+aBeyw2ZAd
G9Rk2TOZdSHBcalULVuefCFnTQbNdF8QwFHqoKcyRIVo1HGvnJCjEvK8T8Wt0wVLYQU0SgIfmPHi
t290LT8smyZntHzzk2/RX+FGeIcVN5kk6AxCVyJya6iHLmeobau8ZNa966ciXve1CFT3Xp+gP5+7
fjQao65F4cneJDr2U2rZ8JvOe7DfBwDsSYhWPIbCGdjJCsNXwtrYhiC40uWrOIfZWAFRlhBL96f1
SHzUSOqzfB4akBUYGuk/tp9XdWJjMvoCdaMdb6U2MkDwuRZ+fnZu1zjZzerTZdTfzcFwudXC1NwU
WMrHta879TIghmXtuQc8lRO3FfIvCWwiqTr+oweXwg6qTzG/cr5IOPdle8ZUEw0Dkc+55kHts3AR
JKVIcOCpf+uJEWgAwnxpADao7rlM9dddW6q4/E+51QIA14I1Gwb8nNp0ZcenzgDzTRvUWNahw8Ux
5taWRDh+WeSMrvRMVdrHcUMTb+nCVk3hmBTE5499mFWICRhlhfwGt5ud1zvzQTkBVqHMuZGGrOEX
50zDlyw/LrHqX1xIf35JJZUGQ5StKy3EdbUYzWPe8rWHtOVkFDg2rcoyx+NbbAMAe73k7sIMsA2w
YgJibXNQmkxtzLJLE1QuQjBgygI5AxCXljZdv6R1hKL0xL43FISu/BM6nGtUpzBkfGvFYrGCBCFP
xtiu+ItxSHaB6LzPZ8nnbpAfYhFioxmxqjQM00WRho8meWZmCtfFr5Gu1bdcmTLYYWe8kiB5P7hx
/OtEusDfvhYP4vF3cld19KeUpBSpa/inTakiLOYkwgyPScqQOlJtYjYDrpi9NxKEasERIO+tdDAg
y7qjCONTn2BMJ+Y47DiuF1NpdpyPWJVkjA2rPcGF3roY1HHmikcHQMP72VONECc0zEn0/BFyxRsP
jPlhNYv45wCqRFyrdl0kbX1maRuJgyF2fA8OBWKyBVsS0wKkDkB7qrudtB/B66bUt/6GtgZ9/1m7
fsjgZks7D/Q/2JAwIhy1EI/TLPUb7jhSyUfTxxarHl0fBY5CA7HGZWerb+3Pw5aDInaL41nxP+LT
YWPqS3OjM2QZ3rWrJyqXuSFnAN7LW/2AHvu3Lgy1H4rjIjrfDyDyoI8HbJqq6gxOVGgC18gb562U
kqLgFBjNo90GlQgqiSinsT7nvvF0pz+RWlBOofWisdwAdob80LWUyXGCi1qND1XZ35RuvKSkJVlt
m/q+0J1gXmJ1xhQ7vsKrkIH/qY7vxWW4/Pqx8Y7DapB2e/bjepzXHCUQHukjOJ5h2O5tTJtAcQXY
BB3EoBRZMB26UQhzQZHGxbqxeQRcJrkUE0HjjKzvrnDS1JyA3KofcFzpXiilH0iBpNelpFyMMohe
ddZboLyq3bRRatAwbjDqB4+WtkCFXZt+H1eOEcQUYL7wenlXJqLszBfc+odiBFd00A5SnDH8sZr2
jDSQfTh3Gd/NenxALdkqITvPg9Hqsx70PV68f528smN336tyfXre2uuU1PTL03A8fUjEr+ncRohY
b8SLMQKP2BdlgB4Vns0uPvM/esx7MkTY779+Va+DLZmiF9wFYQa4JQtRHHFsbFGhYH77pQRtWTXZ
elxv9FEjFgm9GVdqFrqtPAHlClLeP2c3qIxCjK2d9WhkQ2Zb+moFooM3+WBmAhSwjL15qF1ShvK3
OJt0JQ6WCzzzBO2xoO+UK/0iXy0k8T1zSbvcZHnqFQQVYznsZlLefd3G2RNRkee3qUZtnJAEENkX
dkBm1AoLYedHsb2SXY0XXwfvm/jslG+kZCjBXyQJ4VmL0bHEBzEgHxmcK1r7/Jv0oMFHkXeQ00pm
hRShHSz+yBGpaKDCExMU3ucsYPsEsvj8difYgetKddfts94EXDwZP/x3uGjom+WRpvqgNvLaGeRl
en1qgcNiGECsJ5SyobqI1VJnpr47BMlW2bkI5+KlHGed4D4SIUKelZoQCxpSiz4PJxRJPfococz2
PzjOVMMFjP5yRQz8/xI++E9tJz9xO+eOzUhMLFDkZ3/LyXKRkh/it/t1g4DRmvY9hIuGAWXtGWdb
j5mNXiCC8oOwXf7ojAJp0jFkyrZARsbTw328QJO90d3j5CgDvqFqEWDwk1HU+MDJnk8nzV5/shON
jKX88s0B1wFPtvAHBEza5rTc4vqWLEqJGG3IE73zV7Jn9w1HN1S/LcLH6jBqP4Hwu6+Kqd1OTCG+
XssPVBDnL8JAJw1LKjZK0K/I+gPMJY+2xw9ClTQkZ8vxZ8/Lld/j8NLFsl9PEv5G40msNZckr2/j
8tKS0IcKpyYyonUz/H4pLTaYDbQ9BnZy2u9eqQwohOQP5mHhW7N5k03PROwNw0bjRFg/GGlfAoDq
pP6Ry3Mh49mNVcqJ3vAgJ6nVsoggk+stmVoxUpBdiX/kuz74zQvFeHv5bfhUfpzeTpuEHXlUqrKC
NqeXpJNUgoWCdWC7Gthf/RepQA4tICQs7tIKyCv0jnTcYvQoNuLp7l1MYfEGOZ8SnqLgRm6LncJ8
6psqQUH8x61gBg7Afu0rJ4AIpP8QuHzgrFoHnvm6nfxt2t2ttZNqwN+3CCSczVbFd1bDJo18aW+u
ATCDq1FDQhCayjM4lalGQ3IS+dmrLSPOekdnwTjocGzQsoDjUJi9ois/imUTZqK9ccgj0SZyFIKG
Q+uuIHiasIbb936EA/UUtuPOSJxHLjlMa/KKvvdzvDc7qQvU5nTzvw/pDT4D3AFCIJA9cnMcTEBL
UGAw55baHvs1U1iW3KoJ1bwm+/cH7Karq9uAQUDF1uczHxqk2iWUBXs+9aPOFqBihdbV0PjcPLQO
gnjPZuFlu+leM8qLE1vfrWsCHXA5Cfg85bolzH506nCb32jxKaCT2n9w7l+QpRLYKoIEJIFDueZ2
TIjRpD4cnvgz/EXp3d++6zCI3rFkHB52XkyTYJEj3Yp4QpQphYOI6ybhEDsCz7OPMdVGbrriFfJ7
rmEofwlRVwHYGQ397Cj13nr7a1QcZDy6K9jbbkqbxwRxtRNbz6ii2TEOAFlRdwGUAB2DNDcX5OZB
VlNzIu52gseEhTtmMpLTU9ouvsmyNyG3v8qBfVFuH3wlbDSdEK/RgfxPhPg52zpoCEuINhm4fZva
cBYmUtby/lWwJo5gdpqdM553T5hb434Pu7kgskDagEN+hQcZIWZ89J67SGuXgrhC0VayVCsWmEz0
mrtDBpwDvy/fQasykK4HkvowW+p5prlsRIohv6++o2B0g4ZYe6CuMNO8Adg7lrXnNXFCIf3s8Loh
SI6lIRNIYWQUQhypi2vD8BzHisyWrkSDRrJoH92THsdFQvu+KNYPZAU1/4EAljE6yOj7SNep040G
PDBmLmE2INjytN9oo8h/V+kpV/x6eDWbN2tCaEk8wzz8JaWuRvitwA6dtp7SZpqzZ8clkYEUy5/1
g9NOP11dFAhpqezCMLLqiCm6E/7FAzDGv/hALnjHDD+yb5C17eq2ir+d8mNbPLJ2jsDjaZZVUrf9
Cw+MM5UNz/X/u9okgTeukBQqjesPDXdlTo7w0EfrrSG28e/xeOFwxegqo4f097cMtCghHXhsGh7V
C6bNm/sdOLTAefq60rDgvYAt1mGe+pCtZu2yCtaHtIw7EWAwdR7aqGOad8hjSDihAyTPzYvefAA6
PSgoUwt5yPgvZgQi8+YKHWMZAMDWToQsPSUmV0ryt1d1HUjSb7JeK6cBvk1B29HA9gh75Dz5+Xnz
AHhOcpZiaz5z5wqMwr7mIBIobiA51LFbtDu3sn6pEIWv8ls7+dwLhneAzSgwmj1Al1g9CQJV8Qrx
wnSbXgTS8o9qIRiYeriMHTiUY90XS85Ipr2GShngVWKgjn116OlMGG7ZbGimtnk+PM/gYCoHJ7ZY
q1RoSiayWq7ZbUmIFquyGxpgfc1lH24vwTJPn6u7wnYtv8rAsxHxCG5/LSKBUh5wb1osJIMqc+cl
VIlhjUOAyQastTVl16CVO0CUwch7PpxrUyJNOosBsH297z9LGPtK5yq9CP4qKz+acYf89qf6ukVH
r9RHUd8+H6Jb+qM8HZqgQz1vpEBeM9bHzjj1B+A6yR5URSCvZi0hqhKXSNOFLKt1isHWrnK1+R39
rH7xVyfK4dal7yzuZLnfHlehszHIcApkSB+et82MtDnsQ+64wYXFduKGSFAjZEdcadwkdpbzg/v1
EfYvNWJahMvfXLuqKCmHZ3Xr+cpBeFDIesOS9FfXbulDWUTJvpcjI9NUoAZud2kWaLfKTxOfqn/C
DcO9krD5m0QAyqt2wQL8k8P5jph7xZegO3+wEYquUQ79IW2x9MnjlGiodA10qNgEnsNc2ANoCKn+
A0nZ14llF22ga6nPDjfYFjdFnKyNtIy5aNcI3sIReN39GGzOQ1D3/qSvQsHiRiO5PJIHNiH+GNj4
HLYLZq3q9Hu8IiQAZ28LbyPNZoalCYR/tFNLH0HO36+3utOE+jwYTD8v9PALE+lPPlHLqvLpSMpo
kka7AZfBKzKLkY8Y+U/fGPKP83bKGinXqeQ6UcHE2l6ZKLWp5lsArtZROUQ3TXH5fwiUQxWEUzqW
vK+Ky95k+waFIW/bFzjcRbMuFRoIDCPx5kMrMWbeUjBUC88mzekg4NitjG5StA9R46NRdXn/nDZo
oKYLO0oHadjFxSPEgh+2gm0CWNa4MCJGICRoVvAirO0lB/wlaJZ21pvER9lTkgE4mPmeJzrga19e
P5Q6StWDKKn1UEUmHruLY4ORqY1GYA93qdwpNyCvtzzcQo2NDN/tdBTR6aZ0ZajeN00XQapgdMk4
h8rRiLQVe1MGEGIKgq7AVxsMh410/PfYLs+0sKLTkC1MV7qw05Yb4C8NDbCSZiB9JIDxiTzNQ9JN
MG/M86pGMQ1BJdt4nXHrrMhatf3FjzFLntNSKi7ST0sYBptdX5zPkNmMrvlV4FegqVRRmBzCTrXh
nQu+cKUFMyqP3S5P9nP5M+u0vIW1zEyCvB0ZEage1YqCnIi+SkZB2XD0GtdxgzhEqyL1HKh0BXi4
xtvqYw4Srhvv1SKUk65oatbtVhiZqAPfvF0clHAkfRgEIBRagS2usoq4G+ATT/cp5DXMuZKsNUzC
74DisvR+RbtN47yw18NKXghmEN1iFmxsg3ww9i3kFFkthuqLR3afkZkqrzqJsIZHpALeeHfeDZ92
a8CM3bONgU6Je1yHpkd/9BXeRdM/FoRjiCUVRnuWQFKkUaOh3ibTeK94+G1Dl7HOLfOxY/5PgZNU
PT12BNIUkICMQG2QKoCU6oUiOZPHrM2Sembtc8x4v8Piwzv6Rdf2Lq3Zo7WGBetnB6oJ3JeCOZBv
Km9IEaJqp1VBk38Uv3DrNomNJtURSaN3hBt0wNoYdfU8ZXDWUitHlbl7vcS2Y2Jq48pCBdHsvHs1
vsmxDo9Z+TMyoNG+oChPgS8dKcRMMLGBdJSBldCQEBmDKGoD53+9LN3gt7bmlupG8iZsCsw+OiRv
OrLqzulr47xufvnZVBDP2nFkfIZ75eTJDE8zvkDvFbLsnJ8EsbCPR7eWA66kCvsqcU6qsX07BdgW
lk0YoDcGPZ0D70NAajimGmaCy7TCmSWltT+ccsQZLZ4VOMaTb7feQCIgTY2f5OSNHho8z7l2E0jC
Xont++PkKlNwypOz4MI2J9d4PZwqP4iUYTTMsyUr4e0T6OVBOABeVnwU0fnahkVxUJfgOSdDK7+c
5W5Sdfg7xj/QSHGpRtFA/rCa4ck/oL8Hk7CzZM84cRRr3M6/yaIepuvAJipvqI9O+bp2YFxa52Bn
VDZu2kAY9lsv9PxIw8nas+CNYussrCBT/ZpFHD7oRl2mkQIizdZIhJnxfG98Xo59A7cHw7BmIyqD
45ZUmcVbOxif0kk3vG/UALJirjwjfqXRnm3Odt7ewO2QlSJxtvmmRIsm4iebPMp0+xGFGNo1poGB
lqJH0N62Xh3jIynR+ZZVStV0FDKP0nV5aB+9BU6evT5NU+bTfRfDxjjyVVs8Xylmu2TTS1ox7ezr
7HdRutOF9FVVW9WU10yTf0ibbQlSODOoVXBDRljADNCVE7tCdPvMOQvw4NhiaXpW7EAkEo7wC2Kl
NWrGQW0so44nmfd5bJIjwyU6p2iLbTdg+8bsDDb2vc7Z9A4F4t8YiMZHoTfEWlnj5SDRcx5A8wCL
/3DqhCduNa12AQyfzX/Ux+qdT3HPKAYZ/X0KycYF4sg0kQtxLTSTA+g8dt06tzc6eeFg7DiZBgeq
aQyFDjJGCADbGJ2SWtgo93TUUuupCiaCLBqzc6aK7ap07/ougG16W0Pdlk126CYMJV+ML1BThi0H
danUxZ9OwtB8iKJER33LSKMpy3SqyI/XeX7lwP10pnglePKabsN8BkWMfeZswlokwCIaYjx6SCOJ
/0M4UmGVo7w+z0QAXH9SCynqN6pK2Q2ZfxfEepu2zxZ3X42kx1/tNX3MmB9KZ3lJQu1TTv5prLRR
IKme+4Bvxm7OXYe9EoZvRqPShf4cpPPdztina9nSAAX0ZG0OaoRtbNOniYICn0jZGGXaC6XanyOm
TJNHYpOnyrv0mLEeSjOFRZmPJ71bNRBlRkozq5IhYhM3lfoGW5V97c6cNCwRPpPAeejEpjHx0Ivn
Ry2/5+vVbco987UoUpOQwJAzLKdcXnz1QhfPE313Jmtq54zwFxY6Ch/cw/u/y4y6a2g7eJ6OPvvT
LAoOM31rExp6tQlUz/2PZNHOlJExBC2AmItlNKENxbMJhtO2t1KShCBPIrBw4frwgXwc6dBCkNeA
sCVGYSsInInJxsU8lJGUz+gGvZs/YlUTJ+ShlEyrKuoDKvdZ6zieTjfgc3grii7mN7JUexazMxcl
OoWOS95dJrr2bh6qqCUlWp8gQVtBE9kwULtclgrLDam6G5QRKQ0j2ckD8tmoc1JvnfFdNdLBeXeN
BDzqGfJ1XXcWYCSZ4c0zQf1xJDvqT9dppKQ+PI93ErCtMM8AfdRiDP7triNyn/lyQoB/Y9Vb7506
wE9IvZSqh6v5m3aDfkQIN7Uh5vFLu1XYrIeFQAq4i09Y9FZvnlL8gq+4xMEXuIVhlKLqcHjorpQo
g2IVagNMqfcAWgA15pfnDGrWoRz6jppeyOwP17+Piuhr7XcA+Q/o88fisybnHe2iLpZams556mai
eYnvmh2Ay3cH0HAlp8xUOIsF7Z7RJdDi5fRHgirOALYca++zFbixaifsynC1yVVsEFnMOClGlF3j
ocLrxnR+hR5GcBhYFX5YmDLuqS7kjXq1JAqxvwTHsmhIE0gp1tZem2mNPO1nx4VLFzzL8emOI2HR
ziO+G0Hxr00gRUbi5An+6QYf8EOp0ZA2DDV5vRsF8LU8kr2gcfsnquzz1mttkdRhoBe3oAtQNvT6
d4TjmQJmeliuiN02qgk97mNHVE0jHtQxUWYar73GW7xemFeCEejNlDrL3hsxxZiY9UL6MNU+XWB9
ETtAKhcOpOghBt9FkUn1AS85o8BnX51zVEcG2XRMFbRKscRi8//IgoFdzc0iyurbgOfdyOC7U1Yx
tUpM7Gr1zcSVkAfXDgpMOmhOWl+LA4dYaYk9KED4YExMPh0K4WO7hWKWPfC/VoDOWazy/9nVNVNI
de+u06JwiDAppN3hGEYrcMVNrc+sUwPoJu7TXIahwBtiEytpomxdx2u2qV+mSwZbBAq0T6L6qQsd
TDOZQZRRvaLxBX2On9p63KXDYdhsCx24zxJKtPVEqxnrdn2K+HULP+o3qR65UBQF7K0WCG8agi+u
pWiyn+3MUzr75V7cQWfaIaMLOmSs/vDIOYKUN0WEKiyvytqIXQXpAVm0dA+/qw1MhZ9ohZfB3hXZ
w0EO19tc3gAfTlQrdKChdKQUMAeHKiinlksHuLQ9+DW16EqUP0aZu/S++t3tneZv9jw9Xbhyn6o4
FUdLCrHBvox2MezNawqlX9oHSILTHtCFLZA4hNXC0VY4vCp/gaicH3kKpsQyPCWMmkz6ApLDdCxd
pm8lJEOVnyEfR0odGKiKx6yip3RG+h6u+Whb3hc2LuNehedQAESIb/zTI8bpcqQcGoTcAFxiGMfz
agbLWdcW0Bne1/ynK32nxa0xtvMkVBmssfiR03aGKXTKJX7cvH+7dxbikaoLBsLA/6mlqCjIQX+b
q7X5V7Pm/H3ewNUQxKQvadkJYCeOg3mzCk+aT0rZWXDH83CjOUxS4M/MUiGT86npkvUjhV+n/Ejr
qJlWhF1tZQskKxQ0UNnuO/3+mY3oCFKSJxGH46+32SyFKlnLT6tsoyS9u5oRuvOrhGzEIiNALGmn
Z5RsHUstCWqYrwxEeuiGtEPxtNcglhc+20yFPAbi1amYa38e8TeuEfT+6L/z77mxi6Bq8Gm9WEH3
p1+fsE3PDRr/cDcHlLXQ84g7VU/tUjMTLFhibP5IeTHUmAyL1rAPz4wwSsxQ7by60f6RNkfpq9yI
h8OB49TIoF0xH1OvyOGgcnLEYw/arawZ6aDQ3pwp5gauy0mpwE2/QpNoxy0ING5010PnkhW0I3IL
D7oOLkQVytpusXiETi644l+eNKk2ethvJ5WhDbwfJRvV4Svg691EGtgjdrDvDhb0/0W+Ms9P/SwN
XUAZUPvQk8OANoqBN2oKstIMJgP3vsQNHdqWXQsQQCHBjRf/7Rept8KJnm0xDyZ48EbAYCnZvUNM
H9Ay603ryIrgE32YGHP77PcRYh+RsEd2UrJPY5qEuFOo4W7Ox6PTfwxIdEMTYwkUovl105ZFYfPX
tQansjsw3HsoDHUURgaa3i9VEEtfWAQzpBUENMPo9im4YIb0fKUIL9CXVPKJjpxdlYQZrp3nYL/K
nAiKwCd+OxE8b5ZdVdHF75W/sN6todp9acz3nexSVvOAFw/m53MJh3QI2w6KOweXDhK5WTTbwp3c
2+kl6J/bXwdCAicW2uDuqocimM6q+6JlTPXB0vVDIE8oq5MD3dfANJiZK/uO1So7wTJwhOOWmDji
3MA+bBrPWN9zI71qcijWhEW3yx9oO9ayFaqIYJhPoZsXD78rrfDK2NCEKLfwYta3KKB3dn5bUsAK
ptX1h0e5YBJvP4WxFhxGy5go+Qh614AMpXSKK4452sM1os5bH3CvbFPQU1LWPCmF3s2dbHvhjrIM
bHDWcWZQ3mmAHVq5FPA8+0BGdEXkO7XKFDfvdFUNjH0a8iMl/iFEPaV9wUVGISdjTyxoWmbjXbs1
59XlyN+IUVHJ9vyv5MEKguimkRwB7pz8IzUXGgcQ0xnHdTuijykFkMW9wJS4C8xp2nMGkwANjYKb
SEYgtNYVOtA54x9JW7yX8MWdlN0+Tx/N0UhKpun6KenN2cIlFtBWSNVVzeryFsroaPVBbQiMUMyJ
I2aLFIzc8JZeE5q6E1hUCLAibpEQn2gbYM//J2/tI/6DBHuVjTcNFBtWTa0J1yYdowiSPzVooOn2
V1FKSR8DeDNRMVgrgQmje70tNC39jvY65auIp+bCiUTLntPGxRjjamT6WRK2ANU/nkyDlYKzcsTE
VARfd/xIOSr6kWI4VvuGwO9q/DI1Gd1Q6qZdLZqJkR0EzgcachHwNKrTfGoW6204q2F+Xf7rGLvh
QNPGlp7m8tjmiopDTgo7FmrW/lbfJlQgNweQn5vSkX9NO2VrEhk2tj07NXhxTuVlbOfpVemrBpxX
UAVt5E6lD69oS9aPLMGvW4s2qfN1NoeuRfS9EFrwgFS9LK/PC+BC9QH9pjbEmPJNoj2ATSuQ8zLC
XDc0rEsDQhmooCTw5HlZxJslBzwDMKUv5gNQp7xU6oqMaNkTn7Nxx93pv3+d9Mp5PQoKcHzI9q86
w9Q8lgoisX53r8qy8lVA6aGb468YjUHjQwIF0jHbUQSHmgInICi7OVgvCNL259pysCom7LOQw7dU
Y/mWgQuxiRiqJNzbWQiknr+x9sMIRIPvhSozNYvMHnKSeO4YmC/wuoA64ILWm6t6gTjmw6b2fc+k
6v4tvspBkDm2H6Z6qe1NPMZd5KT8k5LRfSMNiRwXRBnyiMR0ak4OZIgb2yRr63b7gnphYLG4mz3a
g1Kl/s1qzDfA5m3y+dmlZRqvsyvuvxKTMEatVFBrXQst0R6fqHemuK3R4p3Y7R1Iw4QUI3MNOCRX
TZjWnurPOMqEx8q/ASxXDqtMwiRKQ8f4lYkmC3iEx4BToyXq6nYlsotS8WgmnCDXKH9R+aHu+IOp
to+6rSTR84HsmLxSh7BurzykEKxWFTmJhTNpTbr5fO7qo6GrRZkMe5oh7RlztYfkfaz/K3TJwSQN
tSIbOtSuq2u6WS8v6wqK3Li5Ocjzi8sN0N+S57Y7qAo1vCGNm0spUG/xXPyo85QmAXqlwLQPPX9/
FDOcezNXzn/pLnn5d9FzlcoxMZrkvlYsxqHh6LyCWa7VZYtegl8Fd6o+Ieo1/fFsN3D3XV7kKZjf
W/Q4OTBXSPOpZlTPaoA8albpbCQU9oySLNf6qvfiAgFzxjeifdNmiA8GGfrPGU4elRFZoypvhOER
b06CpT6jH96sXivAzkMPgKC+KaX0O8shaDP9lTEkKD6kcZ+viSZbByCXTMrxUF38hXCCIlAVdZgd
FmcqMAgHCXt/cKM7FE5pzR6+cJOLHRRBvamOGVocu6zxJGGkTj0VgZO9GIASCYUEqVJg8Ge6wtZI
YhdsfQ6n1+XbyuM/jSrE1nIzDQRwlv/s9Q5yXaY1b8QmGSDpvwLh2ZFjKt7jx71NRiBM9HvCllsH
flg1iu1hU+WOn+hl8meCGtCYT1lvAyhxNU2nXBd/c7thL2KUBlWZW/LYndvZ+pUr8OAXp8hGZTrg
6OT93cRkUbqJDiVBu33lzaCG9FWrMqxEdvzcmTm4p2f8Neg4RIgSl27X8X6nSZH57PHY6L+bu2S4
vYmzx6o+tZ5WYx4QMUwnS0+gua7flng1n2eF4CSBPsc85sfIFZ2gIevs5UWSJ9BV+Cojyj3FxyJK
vs4hQzAUUMM9wsZZsfNxQIeJ3EjlFMeExrUbYbaOA3cuGGB0DZOTWre69NI6/XE/9wbLxSCftIyZ
g8wpjUzej+uTR80mcmHsFj2g6zxQvrptG/t/78zhXNSgeshHpelP9fVARuieOyCMNj7kEAfxINi/
GAPin7xyfds7ytkTBNh5Qg6pihLyMVBbG59IyuIcb8LRSpN1eti+RkhHUOdTVHYk2XiqYF1dCnp/
4Kc7rQtlOQssi3CS9vSVFq1l7Ns5AtF+vLVt/62dBHy807c754WSCt0eWyK8KBKXNf3imcnVR187
R7laCSQfgYl90W73nNXUkE1Q0mvrbnUdE+D/5BINuIjYNHUmREwCyn1EPu+GKAEqPCTVjJ5Au//p
V/5XbSoVHElys2RU373gh2lFUL/rJR3dvRJDBmaT6wis3Y/Ri1sG0nOfrnYpAC2gWRLwgPHd68Ai
HE8yXqI0KxfrVmUAshIeXso0jcKDyxgtPJLxoE9ktYY8UnRRDyGcayOP0wWuEcAb1TcXAhzqlG/8
voCeA1br5eJSO3sqoZPcDA2W5bsBci9IuhAl78XyKN7RtVVTmO3hlneoycH4euUVCztlV1gWeNgx
G2x20CjMBl5hOSMWRHcOU1rzpv1IszZ5XpogoMBvrSM1G8Jn0VYx/JSDXLtgiFc0TSxI/F0Iq1x7
8p3pDzNe/Ig3Pusq0I7CWgTMncMdcfb3Hp2951vCzDO36nT5F3fHSXOpVSnM7fsrjUMK1yYb3vJl
sQkoeU29i3F7gC3MCR5srZmi1Q4VjHXUEEovu5Ckwcq256AvuKgoqFaiBMkEg+8wJYN2bBdsODTB
w3SPjpzGxcpy9WLbDuACwuxy8XI5/hQ/592gD/cqWXGZ303AbucL+pNEaecTItOptGSGBcb6OfyL
T7Lgkc7DkZ776VxRBW8JYDlDXFJxkIpWVOmpZSoAfn85ZuREtb3OaviyXJSicFqpcrxfZ0ujqS4M
CR6BJ0B5TmNtb5Y/MZVfLeyLeaq0257VU5PSZ74B5ph2IWCUIXXv43WZfUjyp0CC6F0ZYXzblm3s
yBRe1FfwVrioU8p5jopTjf5sd++SGjgxf4LQDDpXrPlGFhteuIz9z2bQVAIXMcaObzwD59gUa7zX
GHqPnMOd3eVkJct9YId4ThpHVtxPJ6blOZVMw8LllzqmmdoHZPqKyNHk34Tnro32Mn3NFL9FgXQ1
isYpny/80wxq6Xuw+ST/7k05Ih9J7ImtLKgMWLlsdagiz9vLZJ7XdsP3/k26yOXebYzmSQ5Ee59V
ZCsILu4YQh0jZ3ItWcLbpomqF7H7PK5DCRP3WNHhL8y0RAsqg/huEIOVaTGgXHyLJfMtntLt4Rq4
NoojVZmY27qlx2i8qVMP61/AJbSHSuDUlPuafMoJUWfSpuSl2ZxQUURzcbDDjbeCiGInJ5tMEZQS
tNLHvcGOeNxxfKFyeNz0l6WZ4IeFHPmHa6C9kpZGhjO0X5NzUByPw4gudl+TwfvUt3EK22+InipY
JuT4OAeCQ5/O1j0r7AiQJjGFPIAib2UWKd7X8CBnVtaZL3HFE9OaN8SVAaDD7SxUE/GEjESLG2Ep
p37BeVJBScb/AlTilxYrvJxF5fSdo5VnUhRKFgtHqA46DUO5AG3XhBhiyp1NiSeGBcW3cZcsT+l/
bnUaHkQFLwSeVzTj+JYimt7f5jNEoDrDQ2Vj1QtxD6KR5OOrXuUVH+RWKTLSpQ8L9h2cUml/TkdJ
mgU1GumdNg2d/ZWY9EQ5I80EpkenBCQaxH4HX7jN2wV6diW+yfu4yF+pb0iUv3TpRFjNd+Fm2S5J
ZSsiXOI4sa7DZdamT4Wan7W4lrEzErVEllgnJfSZf08i4EK+Z+Xr+66ZJ0Lq2SuzL3T05b/FAQXI
7x9O17X3maM6tU/boIFYX9ooAk0JwKrARoPFUoKZV2dsHrXBK2zfsa2d/8JzUMLZ20zzVTsXXM0Q
V4mUL4/j7kQ6T1BYmgq1qPS76vNufY7OBSAywBK1+sWV/7bvDtuK+uwgg+o0HnWmUdSmBr4CVcaR
RiRT7b446J1/tppgpZov9PS9jRZxbNQXe0ous/7CBnt372KxsAfwWH7WbfIV+lmBC/Fw/TDfWAQl
Mzzg4iuufGQBqFfibm0wVecrNHlT3BVGDQS1GC2jmUp2TFBHufxvJrcKOLdpPNlXxe/wop/aSSpy
awAoa6QY4MJ7DNis9PFifuVj//dLX+ZhLCzPQITXVrnBaqhoSwLM0vN80nsXoDlyoMh1UF/Xi30D
7s6uKHhvroqQ+KYvGyP+UAx3DFJewiTUbdWt3DMjmMcKJN5nBRcbO93ADPAgbkdtQ52rUJV5tq4u
i5AYVqV4ovG894uNKhZ5L/9IOV3EBSMTggea/2gnBVFr1C9v6i4VapQ0cjFMUyWdktTLvU6eI53Q
vOTsI06n+DSdtdOH8P6JXRKPJ1e4PAj5QjZFHWb95L8zwyJO8OK0SRtfnGV5KCtQY5vYaF+1eMJn
BpXE4PJ4Y90P97hO0RvCTsyCywaG0pTlZqOKvA930sEoXbO6GpY6otfDDQ2BqmKBQdJ+2Moj9L3D
qluwupIhNhg83drelLI9Ck+bjhgeaMt6JGBs+MQgNDVxgNkDb+WbNxEAl2WW6C+Cuu6+K53gse9i
+b755Sy86uUm87qH8bDQtOcc3098gubx4GPhH5J8PItc/zoINstYqRrQvGI2cR8Vi2FTQE0t3bho
EHxcqFT+TnJEtksZWXggeCqsRYpgXFRsTzFDS2HaDlHPDmud1q/FjTLZfFZCs0bZxC7o0p8QW71A
Ql/KiXCxCML+ZSdU8WtVHU2LBTJtzruCW217y5DW+kkcfNpYD/wW852UXcFlcx3NAVS9968cZOaD
XjOgEj3ARSiU85xylmZlYOxRW0d4JBZ6M/TEsV/QHwfp/Ue3/zpWFPmyhJQ5XFzlP+/7FAxkLv6M
jrhboeJQpgl1/rtl48Hvvm1Q+ACcYHrzTbjRnyOaxWbVVEwE+G0/56moLgHVJO64g9NTa3J3v/40
4ghwHtOGsxWvGso6VRJk4UvempkfqE3mmKfBVf5kChPfH6/hZ8+crOdgwJr+jzSWRFRDTPmfXYBa
EjT3R0DQJwXGDlItm8lUD5GVhQAX1L+wJdaiJNbBb95QL6ikb8Ho+GlPNkE/lwbYAFmI0L8r7GkV
3rcWICLsHGeANAp7KrWRU3tpgpsKqzCm/l1FwIxaND46Hd0gxdJIMWVkIewf7wP6s3ierrIiLvI8
Y6l6H69Lod1KgkYlwpLvEE+8avdNjIrICxBULuKV5vWU4w1oxFDhj62mw2GxaI8NySP2H+DDZKsG
E5xipkHA6l1H+VTC93YrL/p/O9aIUdRRzWML3RD16Gm//+jbQWEg4WXfBPtl+xZL3fbI3C7yQQIa
47UnCLDNMKsk1BNiwM4W9mDFU8Gin9Ka79rM43s/iVc4nLkta9OrdpgFh24z8PLJLhE74LagS4Fx
nhNNq9Emvig20I5hpWHSEp3lwS143ZHgA1M0bdk7W1V1Ic1AeRSk8ohsHBLh5/50S3CS+r7l/u9v
LIRndLUmdCL6y2rGN2U1oYlNdYt9b59F88oYwJwOADxB9vKeq9Qp3UhZVKTLH7qdbL8Y8whXzUDN
8YB8U5M3YFscwNg8m1ciuMA7sB+x2A8ayr3N3dFx0Swc+srWJ6wJS0GrqAWPl9L1N4seJ+cb1CGe
i5KNEFKk2XpGyv9d2gXXQGasVBKgDUYInkhetWkbIitbotrxP43+0y9TTZR8599ArZ9jIh3FznAA
QHIVvsDr6IXL1Ln4JPFAmqCs0P6JR9hnGdY7V7uEE/hNZKCd+TnmFTLTL1X8KLjj1MFeUX5EwsR5
04wbN9p9Ggp7e5pAixLklycB6BMnSIFdPTCP5vnzqsVMi2zpKIyq25Hz8B0OLX5/D8nnzK4BjMpU
cNoBZ2sopp8IlSY6FE75Xg7ELyl7omLlcskZG3z0lMTr34FnYk6nPbB1zMdg/GQ2yZJY0BIeuBcN
PvU5/6EDiWkNclmG822c2DTUyJRMKywVSej3z7vsvYe1izbqolQ8pwb1U9FHq5tGYwNvULdqVezx
gngUkcMr3wwFvpnjPz8q2EUoY2vBlsKfxdeAphHjzalyvzlsSIwt8E8qa4Opw9rqti3Yfn4jFSEh
1tvzXEoFe1GHwNKfzuHbHoR0vWO+GE4fGL4ysmZQsHu6CCLsxAlsmpVhy5TmTKLfWPh7Kj9e8ALF
9Uw/TWqr9t2qin82cZD+2AA/ew7Zv0Wzo7vS+L25Rhim6XOAIyHM8CjK6Vk6+CmHRjs/yBWgDudo
w2QoUot8a07+9286tEHIdN9TRlYywh4P/rUOMLf++MO/7XgeUqse1Lf/FgUaADFMpH0Uk4Wq3nng
FynyPIxEOdX9cAfb+jwgp5KtHD1AWQlg3foutRvM3USDkPGVtPEbz467hqE1cNhThKpq+0DipAZP
Bx7paKW1lN9e0QE+rLJD5ldH4vDIZcm2q3ha5ssDn8E99XgSoSow3bbIDdbKgEb6FTCszdyt5PS6
VrV10Jmqi6gqHuqJUmvszpNqTl2CW7atMfhYCMLHkaQTDnkgGVrl3K+4aeet1DHpo1gAhqlbV/6A
rAllFoy5TbyhkcJR6gyqQO3YRN4zQg6eir9DPpKeDLcpizJjcR6FWBNz/R/NERVoNmJbF3y4gntc
eF9AmD0IkFEVvsg50S2P49cxYQfUuPOy8dHS083dik9OR9GRenbe3bIjcCktuYGKX/3CJOpBefda
3xdTiU6oNya2gqU3vctskfn/URNjYalG7C368H4YZFr+LqJB5PW3+2KcERsuFF9Tnfx5IBU0Raig
PvrOaM6MasLWfz1U1/xNfxVCiDRMKQ+2lEqjJD25uVfy7ZIG7wr6TLt905AyP+Ynjhn1ZxvuKJXG
eNzqQTHvhAOd+i+TwX72fSaZ2WCDWV6TEuZ4Uc3YVUzD53GNJdfh9ppGQ/0uI4Smw3jKalDOftYr
zLD1zL4cCOHZlLdXTs6MmK57A9OFnLb6EXaIB+qczp0PsNsxcxnbHSTqrv5Nqn01elNn3ttctlN9
jSvDkDLaRC3pq3/jbgsD5cXl0CmW/ncUCmxeRtc1xod0ghLzBKpIIrbphY5fOay9zIsxA4lVMOLo
Jrkkpw7Zar4RWX8ONMKyE/ea91mq5bQG9pmFE3Uw0Ut9NSCikRtZGdVr1/WnQ1p5x22L4MiD2ZZE
r5862WxKEfJGpv498JOH92oNGblGbQM6hCCMiKXJw0Jbzy6+QziDbIgH9UeN0OwwuMCXGc9FWTyh
B7zgSJw3UamhFF0XYO3bz/NhPAQnBOalh2NK+XWHFUcdFmQMkX1VqkQ8/Lz7id+j1tYjoF3l/TgU
TPrn6he49UedjC86EiWn7+G6ahYd27VHQUso8e15JuCRjoPfW581anDwh+pF2XvuXwyTNONg5ZPz
JdYaRc9JL5mz9F532vVzNDDBwDG53HGYxoPmr9BmeuYBVes5vFhtt05bpeMR7sCAtploSmiIFHzl
dq9fxgPGdoUv35dTp2kMcMN3EbtD4wXYDML2JO/j+41zF6ssmDTM6WCF5Be7/ejnAguuPl8yokWa
BkXn91XB4MRNtEw3H+XooqNhJXTfgLTWTsa3w7KJU51XtDkcLYh8YENhSSKscKXv8uZ6pPagB66o
hpRR0bPLLCZWnm0o96jjp/rXP29smg8TbSEy8or+admbBwT/cith9SnOroOFgUOtdkVm/uSsR1iN
VPH+7GG9X+WIqoW0LKPPoWrx33Fwz87q8E32E+f0hN6+18/GBoLUoIG8qDztMVynVxIXTMBWXpXK
PPs3mFimTVJKwyZ7Utm/mJicrjTcGHu9L96ofOjBawuYu/gV49UxYXGAAVqmCnpdZeG4or8cEzco
2Di3eJ8VdzT69dHb+guY/wZoWb5s5DI0M20ntAweB0Y/aDxCE8fflaL37BsSaHfs4Xa3WaMVP03M
NGm3yK+euHyvUovhSzbz/kxqLPiQ8DomJcxNwwlOcXc0LSQ5jm+vwx8xoHpYMpyaNxgIxKifORnO
ghYQteH1xEzsmjFChnyydSEUe/OvDjfLqpl/XXatJrEMwm1U3hDBcyAT7kTGBkXd7BGfgKiL1+U3
fKF9c8xZNRaLE8zKmU2wtSJp+CqMyj6zbZKPfqb+Ul+gJi7bebOOQ0ddgN+DxVxMNDGeM5tqJjBY
4G/g3M9twCNYZaDzeg/3Un0qdAuFQnCkpK2F3TW3HuliWYtDSvZ1yYXjkpvU8QvSSuh6HsQpYQir
Kk6xe6eOis0EgUpvM6zcMtqXp2su4e6iv4r22uX+7O7NKLkSJSuKM/I7gvZQbqzVDLLlatkdK4Js
5tJ0jPVfNfO9IA3KKP4zJ/VWqczdjCEMNDS5OxgpWDxIoefQEKWGRacs9AwQMTO5lS4ECfHz2DMw
HeyWoC6ID2VOd1zTP2kHmQO/f2PdHGAO8HTsQ9th8odeclNjpXEFR/BzELbKmGcTlOg8snJ0oEyN
tJdxAKV0uahvUW8XphLxhQh44BEQZri3DHTn3Vmi1v+qYwBz23RyiRQZlVToNQWVoR4Jd7vAV7EO
q8Qv2H1ctEBxkBxSZTGGl+jBkSGWugQX4UOyrCK7LFSlopUHV2c3aYo0hkVSh5kkY3PdRZ9oVmw8
8j1n8gb2+A7xRZ1DsuShL4vv4f5nDEZh6FqOwbIusAG+P9kE9YOqSP44O9X8l9sqvf54HyutOL5y
zFwWY17t9F7RwVlYj1VN1zo0GaJrr5ueoEQLEX+SydKgfb0bNdeUdJdJ2U/zXiR0pBVIRB0j1lS5
AKXu1pnsHPQlwaqXniIVGMRggyM0JiI2NMKu/N2WBXfFj7pmj+6NjW0ims5691PJa91HkzEVrtE8
GizqTAwYK7EaPzF2IvueNILuL1M+XPRURNLpQyLolvthhWErldu/6/Gla7rkZtmEkqTbtWm0GKV1
LI21F/jzYI1j0z2VnYX3r74HaPtJAd0jGkpLfcWBs68CGdSZMmlq5HVK/co41ZZxJXkzLFT6u1OU
dncTTc5LoxBbzsyzwj2YsoWeQHql2c8RZJT++L+WnKBIBfJXeE+zjc5CIi+g7LqjvlYnaG4U1O2b
YGMHA4m7J7LTM53xBVItuBbBdjHyEu0UY+63SRNvoN8ilKGMTuTZWRSz/lVbztqMZRt08XfGoxMt
IvA7yCJPgvkW4iZFaETahnVpUulYhqXLn3LLoTmbPwBECcT4dXmb/tDUT2msFA0gcku5PpgQLSdw
7YE08KWFdXSzKVv92szx2Jx4WfPZ7HhRNrZXLCBsPEJhTdUwB/0NWdMF5f1fJJ4tWe2OB1IvVseZ
HGb6eovtpB7fXtB1ylM2jzfhCzL6yWGTe9NELjhbEcbK3ix2QCT2W1as2Dbp/GtCs1EqKBtpmzyb
mjAIwdfSHCQllcX3sdlNbZ0ZfyjaKTGqncTCskQ9+POHYOCamUCQ/dR+DSCbYXUnOfXJKPcgrkw6
jy3O3cOv5r1diZueGtWNnf6Qym/DDM4D53CyZoMe1+IT8FWIPp/6eRf7YTanezQVoxehdM3CMTBW
nZNVR2A69SesaO8wLnXUL4MYch7rP45LlXKCocJklRIBZxETFbv6+wZEonBA138KFFTku4qIT+Yg
nVjyjoFIJT3DAObxTc7re2ZBVLJLlYrh1FZTj9kyB5KIVtioIvrbv3Gyz1ElCOCTlnJ5ggov4VJT
QZhBa3KsRPsEuuSzM8r1L8gAB3em9qbYOgksOqJn/IK424GowoRe7ajnRFCk5cK/R3GyE9FGoW9D
LIYBf5m29cHjDhv3VxnyU900v4a3gY5RNXTD0U4BHjqdwkXpaq3Vg8GSUmMQZwVn8+7YG3FKpUOF
BUluUFqA6wyukiO7vVTo5U6MDprGVxBpfc/BLCxltw7FndRz6OyKOyeb2dtlLSO+Tpc8wO/Zz8R2
QNpvdtXbmpSBBunH7op3DgQicCokTdh21MJCutRwEr7hlOA3d36Wt4mlFXVqqlDtZEFfgPlr5bkX
zJapCoiV2hxSt8J9VCubqNmzTSQK7Dkz4a3D0/72wU/scv6FfUe6xeW8pIRoAZKGw93fJwws3w5I
/1NJ8ceeCPwCTZ4bq5nbj030FDozvrcRugjsBXJBDHc/85TuwA6J0iVgU2Q91oPWZbmLRStez5W1
CeIVnWUX1uG0eJvJTZp+cMs52/McV5x0hh16A3yb+LGEUdTdigv9HLG2QVxE3RDmW9Mqe86FpAPR
7fwZwilJoxocsxKlOW5xQa8+jDqQcZAGJKkPpAYL/kOlIMUDCnaoo1lXO95BGUbISRd48SgD3B+j
tTM7knp/5uj5SPVR0QuzaNEFHgffmM48jQTOZvKv21CHoMCxut6aATBFsRsrOc1Sn3F+W4765PRc
+B0oK8hBz4v0UjvvQ0G07SPjCdiJWCtyWIC3x4Em5ZW+lZyhKQ9iA4vnccaOGgJSNY1JL4OUoAK8
lzKoVJYyQChpQsZa7b++YjYSEEpigKIVMMbBuDhy3xoMRW2o5GFN3qEBMYtsADcQ7tRXNvN/jlJ8
TIY8zwr3DXlIYKcoYF38k+r2OpW2qs0vWvwzjSc/Jc8NQOByRPYVgN0kW1kdPFqFu+KMwyLdyShX
eMBPETjXircf0icCoDyyotcXZTosmesYOvf75E0pSrsajlvFVpdXd3PpIj/O+Yt9kzvpExL6Vrv1
Gux9UAwWKqUsiaGuK1zNBRX97NB3/mpuxdalJtrj5FDQ6ivuXaaR0aeMnw8UJQCAglSK4tnx5toX
CvO3r1150V6aBLeL1BhiG1eymkFa84cdZ2A+C+JNlcx3ERfM75ZzgGNRtUbKQxVdfmi4HpNrnKyu
3hctYJsolRj3EIgShQkTaBkUJwVMAYqSipeuadD9FV4nGS6JAm2T9YdCTAAtG3Mhrl/EFpzcG0e3
J5KrE+vAbwrxamduLga/BVH4StPAS5avQnJhdkfAy+2fjfr4XCgbpg3CxShGtSr8NCt42YTY3bEx
6BNVkyr7jOSMu1YYr1VHSb+afVO80qspBc/OoCEfDoIO6XfPMjKJDp+rpvO+LrXSGudgRsZ7jrIz
l2SqULf74Q8koD7xtCVpZifqz90YK3eTcB1NjMKjkP3vNzzmNIHuNmTAOLeOCJW1m4Z27ESWMdzS
CsuaUzeTGwZ8O00np/sMhnDwpJY6geJah8fbx4G6YM01AcixJyqP8LchOcy04p09qLYKRp84Gc+D
A0ItoaKIwk8DBmDW8JYt6X/gPCRMcRexEAgPmkB5m1/NYHfLVEODm7qrBMF8nQ+hFVnLfLtOURX8
IaybKy/mtOY1nenHYpoq6/bNcjLcNU1uGatTSUBCU5GWILV/uOS+emK8z9E1Bhb7kqZKEVfRvF9V
nls864C8oc9aPbee/RRHhtKpxNrKnKlOECVaBrpK9znZRqwKQJd0oj1u9RpgnF4cdZxJbbRbSdtQ
2ThyU1QxUhDeFBtax5qFHMUY+kuECD5sC+IhHzc7i9SSwcG55yq5cgNyjsoA0+LsporaBjlJFoas
g75tZwu6ZK2P5Y+tJJJRKZVQ5XJALgo5RG8mNZz/L66m80fLgWVJ2WvwZbUw5qZXYBwDOBGpqIUd
yoK0PBmv5dGcCAmhdmV5c8ze7Li0lpycw2hMVZwQDHEg9NusfCIPjxnO2Z/1cfK+sPrbyc/nZEmc
iDTzH6G3uRYTCL8AaWCjCCLLpAFK/MDqCSEVYBYetPQ5ou3SAKe9q2b4rNWlrN0nm5LrCcTrty6O
M/Gj9v/CjhfhHx5/NRpJzHoETP/EOZ0SRbyyrSStOCHyXhciRSDqdRbWwVdbyE3xFblThhkbZr1/
zt4Gbc6IoE5Y7JlBCAjuwwaXd8AeVKqWuZad0cVZ99riSY7L1+nrAM1yuHE7ilCi+eeKVig7zIxD
1QZ+xBXPVscYmUgW2uvNGC+mQFIQ6wrWONWcRVszgqX3noiQcy4RhqVV/FkT2MXDaOL0uYEP3hME
g5yS/OIpDdnNYjUls1mNMYnZNeaMBUh/I4o9oxmH+89Gjt2Dih3410OFpumqUb/Ube4XKFrpfgsq
x/bpMWjLFLijxgBTfbxqtB6vjm4vHXuvxuU85b8LUP1ArVn+9vX1U8P4hEekLB5wz7w3Jo5BAUf4
HP3b5UiY6Spm4jtUy0YH6g4+sBT9iUbuHpHSPU7pt7dYmPW1LdhE9jBD2KmeSLraYenJwIQddwIH
4fBUkhOZ6udtEh1H+3LQSCtERr6bPLqo7Zf7UqZ0BjMUZ0lV63R9G8/n8ARzFIqbb0yAA6UKwQ2Q
ekfKkRvF0qm/6uFkGVZowKlp2vqV6oQ3iRprOQMJPuvJXV9mEeAfN3DhRUqAukJaEBKUN/z+wuwB
jMTy5yEk/OZUplwyy8UDnm0ivEtosX+GjTC9XECTpVIzVyAwQ7p2RV4QvBbYWWmAjGYMABsmqFiO
DrvZORF+BbLlNf001Co3Q4hvmwFBolO6QzGEi2o9pVK1UJyz8tk08mnNW3qk2uyqTa34A5WXC151
coWobkFkwA+X4VFEgDHDyEUyW24Wl3KXWRIgEsWGxGX+wRwmW2RQlDKeuQU4xLy3aNkBjXl6W5dD
uPFHT8ZO7HGJZfAtJCd+7a8ZUGcafSjBeCJSzpW4cO4x+nMgQVMVlzrw5/e6DXl1IJUkYaXvJXBu
j4FWPj2JczJL5c3HZo81b4DsUbMnzEdnGllSRX7IsXbRU5MwZrCH8XdKHabpfa1u9KygAQ36Z0jn
BazCZJ9c9U6KUCrAbjJTIeFEcBWXrzqC93gCcZx1M5RQHtwHodaeRW1zkBuVTH38R3zATaJhHcuK
VZzH6ZbbwNUoFIdVNMij6h2w/9B4K//Jl6mhi5VXmLQlD5g401txCIHf2bgRkfUB0S/Y2IfaluCK
tpJ/t4SatEsKOgnDWbncMf9XAgJrtAyAgEzVX6sGP51pyv3xFFeoIGKptrXT6TwSRitgweQsZnvI
ROqsw/qFHZ83NAnZkrp24xOcFfc9vMTWpP8DGHBb7CGoZ/y00SASCtqc641oEp9/FvADaRv/5ht0
11Hq8hbM/Tkc/BUm1AT+98kyR3BxNelygmwOTUnBMO/wt30SsPql8uTp9ccqGxB9Pw4KZTedEJ6z
oooQ7bmD2W4NzZ13FrxVUPle2Axh8ZJ2MP+anrONKdj20tCW6nwWH5Sr8ruyTEbONrBe96TFX6aP
StR0nFj8LTgM59/gJaNoYUgFJoxuMtOup3wP+rYx4D/Mko/+V9+hgccRLRrZ0WI6aQwzac+pIpC+
o9FdlAEoS4TfPYGnV0f2fY/g0vGqX67q1P6wDrg2azKvCdxLfXW3qlD39XXxSJfyTanBfVWBEBXw
SCHC/qCR/edqSTc0RmESLVsvz0rIE9p4xZkfbD4uXSVB4gbfROjkLRJPOR0EjJsR1QdDv/KYwVS9
AWcaLyCC6N4ECCSvql9uXBMQV3ec1nzUBsGZZGV1G+qO+gYuKlAcFd1z8deybocaC9HWZcoIuURa
/vW3lAP9p5meVbs49Mjw20e1dEN0pYiV4kAvZ7F44I3nCjjeBtdCwIY+6ZpPqXSojCJ9EN5/adKW
sf1vpuBqbfuvo7y4rAsqujkjYpHW6HEebXPqK4di9vvlSXfigleXRL4r8WVtT4/DGP3E5k/G6+R5
LoSiHPIXve0m5Qlx3RAnPxAQtGh5SR2P7AAfiL1PiBOiAAtK846sBGLKAhRCZhyM2VRlPDat9ayr
E74F1DbgLyBp03J7nZ7jlpLVv0XIZ7/ljONZJO3Iti7VZfSYUdpGMvbIaeAKu7B9ptNsbesn9n3y
3DKmxUii4rIKlxziILFkD3q/tX3Tquy9OKrZcjEbgEFVXyq8/1m4zqAjXsf84EZv40vIUhiMLtKG
VKbRCgwL9cu0sl0WuaqP/qRCpabnhxhiaFiXOw3Jh4Ns8VCJNB7nd7Q7eTI6wDuOJGCqIs1GpceX
4t6GpKWbSTfD/2k9BV79eSqA6xW1vO9v+0aN4+EVsNLsejrEv0h3KdPwms0z1rvVXC9TbtaCv85T
qYyPWHm6FCIARQeZdNaPGsQPs6ObSCrnDq8+TNOcVimIyYU4/TIBA/QTmxC8sn5uwRNiZ4BlBXvA
aa+EryIViAe2qULsu0V8zAOZ1qXe2AAWJhFSVFjWuPt/FczkDsSo1oTJrQ+zQnRkj6pEslOXNUeF
CL+rWNABL3CkFkQHhVqq2on4FtxYEux2a7y+jVWsE05YP/t8BMuHOjvzhO0+FDS9LqYeKpY0qLd/
W3dWeLzwV+0eT7ThNqBgs9oKIqdCr8MKU+6uzpdDlMyfE0nlizthAk4lRPHAK/5A6SLvxXFDqHbC
GqC2S7cGopxm8qS1Citc3dvoOULFhU7BnQhY31W0miezQ7bX/bwdr3tQ3nKKFEK8FahRXiBjhAhE
r6qboV9F5+DYNWxjKSIYth5d96z/OvLXqsESjZS/5tk8gWMbcAIvYbyvJOXtK8/y8jtEesViWjag
OdfjFsTrmrcTOVoBqPTdXBfYUypxUCItU8iZRs9Yc9S6PLO0ulW4a/lDRU6i6xNs1I9mckepJ2wd
hh762rQNIX3OQ4tuq3znbBkzRIZZbOq4NaeCCRMZ9uvt2N2C9B1WeYXVkcg4QXWDPZ2yqkVIQ58a
6rAm2h0b8wnUcBBqyuoER9okv0Yqjjh/cs7YwIyWwVWF8fVoUvYZ1mqANaGWeyqdQbdJbNQh1ncK
+kU5GL3h+mt34snz0fAUD5l631CeUVSqq4edVX/LZEdcGD26d0aYSOTKc3uW9G9maAsnwiyhpTWh
XBEYQcIwEMPW+MuUAlgcRKHxTYErzXdHy/7YJ5ILVQE518vl+vHgefG/VKAPGJnII52ufEp2jMGq
DmhuDpSLMGhKAzl36L0WUU42+L8HK12Oc4kz3UOpdQveVyxLgtHVkRkF3LZQ785T391EZm0l24kn
qFR6CET4U16tg0eYzCCTIyLpM68RLyvZ3HIKesDmYbZ0XUeGuLqFg/8/Di5bx4GrcMoafZ76ZEj5
LHajzzf6DDYqotXEAJXfNikC3VYUwc0JDg3mHL6t6kjK8vPcLQ9NemS3TYe0eTGvNndtl6E8wm+z
fCjDyDKaPDbpPGyRvjiO1JFE0xPzC1cnfX5G4Y8MaL8DVzBiti5hcmWfUDB9ZfJcThFPxojTXeZc
0avBhW+9tH4yN9cILb+iYjwqJTn22esDdy+Vu0+zbH16ZDhe64FQ4O1QWpbvBulIwQOuoWYu/m/K
XUlvQCFnbLLKgQ8eu256yfHqTGPSqa7mXZMxhRMZxh57GE6S4oq9yzyJHeQbQIzii2h72dcQIsdh
Qss2EQc3ny3VaS8MY9whnyHMv5/ypK+pq54o3u17mBPhuOw25SMM+JKAYprJEtx5qMbrhVQ9f7fN
wHw6fOgE5uxxcxMRLPWkozPAp41VO9JkApqM39xaJOxjDeeNKKzeMPP7MmaJE51XZ+bkPSy+rfcj
4ttJ1oWTiUXR9r6vR0VF0OmnlrRj/vVTGRZ8Yz7vzSkdROWO37ZwOjg+O1yq1zdHydWmUcFLtAc+
d0Mcwjrrl/ZBepsuPh+y21urw5KlA6OSLv21m23L5Sg0bgLMUENhWVIui0ZFZSfaC/C2lqalO3/4
LYtCw+EML2SlAeZ13VhrxQhvgMjJkzhoqkAY4zhzlxnG0MMawXuqiCV9mT9Jl+KkpZOuz5OgWlcK
34Fi4MsMWVeCuZrRj9GmwoTQRZUGFkfcf/yrTZF2n72YE92cmkB3btkCzJq7UCAsopcgt1zcew0d
Zn5I95befpYajut9M5gz3Nipdp8sA3iQT8JcnkecdafQPsLqqsm25yLyOJ94OMphimOlXXJvzcvI
b0rIdIQMCupgY00gRy+6W+87N87jTnKl+s4bngAc2LQuqvw88V4fVHHI7CLB9/HE4U1aswTnMs10
KOZ8T2V4bR9zOu/cQqD6W3r738YjSj8oSQ0+xvcjO2lPNyIj6ay3/0jTd9RMzLlKekLSYV4yCPro
lsUF5pvcIwBWGmUDIerFAAev5mJENjeGx5Q6OsCmB1k4J9zibt1Hug9Saqx+ECuHJnfrZpDAayI8
48AJ85yR+nsLHx85mzSwRKdqMHH8NB+EFpx+CUTqZduA7NYsVltD72ECMaOrcF3tbw4D0m+V7p6W
dMJIvT/QYP94ZVgBd8e7t7uQ0ncT8+KIHpO8gAunE892KnntBDJrIAQb9wHXogxU65iLO+CsWaNf
KE1QQEOssTb8tBQzuy6MUB+EfWKfUFEjh32yH7mWaswhpTFnyyCm3byin5qqv+xERWD6SgNLKyfF
MN1XhEw8KUy3i2rzLOnSFrRmO2qC8Z/4KGuBztIZZiLq+pVgBX+64Wy+w4qF+fXsoXOmsmJQDDdN
E9MMkqb84IA+LH2HfT8D3gzvVjyxUJuKR+uyQhUJLrda2zMauwQfnKMZwA1WX7UfYrAQ3efVHpW+
bnlMd5hkMQ0hPNK8EWX8H4j+ZL0EdtzBlYjJx/5Ia6swt7pWM9tGdLBr4+XaEEawfNGlBRIx33hY
b01UX8oFSHMm9tS2ghENCDlmcXkzwwBfZq/wITgjqughl65XRAZpiMEL3Yen+r8mLXguPQKh4vMV
4RJQ6xM3GtmmVnWAjAE2y5SkplF4YKTgv9ltjl504QmYAARcfUfwSwpqO2stCMxaBvBch8OMa68K
FilPQSONH8ZatfPGmlwtK224VE/EUN4rg96qPNnBx3iF8rPjddc2B/ZH5Q7rmtiAmhPJU/0pMoNH
4rERZDlkI/wY3gN2SY2nD6dvZf4Jz18S4eEOnTiKnOEol6Oohrh+kP5LibrcmVL3+RlFSYYLJvu4
qVCV//QvII4EKXBGqmeixXeEcYwrQs0TnddYf9vtQdYOkcuwvBahSZ0z5G0iQjKgOVm+vPn3+it2
A4zESxWlOIvxf3lQNiOCp7aWt5CbHGR218+gERZ7zJmbLNPmS0/6SWF21r3zhUqBRvdd7Mwy1UIP
TE8WbNzwZfXxbEDOqLKY0IYQ5ksvY+uXwY2rrYu+YngXXSOv9bBk2IFISwlISaquCk9R1r/pwt/n
8UOnTP9m1ghXw32h45yrNLZIROrWqUxwvKxZy5Rs4FcdtvpeLZNP3INQGBRLV7GDAcCya/4r5ELq
fAuBjla/LPwLM8XtjBnKlUV+UbeKddue4me7hlA2nJPwncSCiZktTa2aKB/rpE1KFjASl/LEwa4E
FQcyETcp44GayDfMLvIRkBXPfbyD1DoHMbmk3VO/gPRLGAU9gFUE+Fa6T9pGZp7v+cxjaTNGeiH1
f12kX6VSyFbT2QXa4KUR4zyklxfr59S6l/A59YwnfOwf+ETmCTx/0ot7NY+S/OgJj72U8gPN4jFI
aodppL4Iu+ElP+pi2kouycDZmhDsvQhoLui0B58t+bSISbSMLyuC5TkLEoXZxhIvVh0p1Ey8ht14
BW26GtVQ1PNLk9yTXIlSxbfrSM59vZSe/d+luGUeRwLtuW3PmqErj701o1JQuVQieVZmBKelUCdo
sBkpgRFqPrvsO1RZuEBkLOx9hgrR3cYfMbJQsIcdsGZTpjl2p4J/qaidjytb6pkFlrTJ2oxj6Cm3
ubk8Jj6qHKLX/8KyzX3EHBehP55pg5z2VH+2gqDNHE2gc36fL1xJ93eBWiYtr1J40mKDG46Jk+WU
GGIgkftl6IylFBfUqyOI7CXFseR0aGWvaKjCRWmrAoXyinJlyi6ba2LkD6crL8/OJPlAFD/rigZd
6uafiThCk7NLnTG70OBVjOPtbW07vmii372RWO5EKIoPzNBKoyIJxe/UgSyx1tAglAJfqWASuJ99
+nqr0kdL6s4VRgoNvIXQegbkF6DsoLVieYERuHsmnb1+hBoFe/MyifrxqeG1RQqQ4SMFUWBuW5sS
fyeai/MZ42iO5NqQnjpn5fCwKVD2dNcgRKI2vwDL2zZHBz2jSJKHBqjUfBKc6ZAcpCyqD55rOCFO
myPTZaVcPKCv4GU+bZykmC6BJVx7or8fYHakJp47e/B7PEPJMm/hCVUXayxRE8azUuylyg4WBKXs
CW+myx0kRQYFzBtZPBHkA2eyS+22CAlu3r/scw7KMXG5RqfvcWBkBMXaM7RUfNaG4zgQhjpECsek
bj9LHrwiI4NjO3eAfdUiGM9+lW5oEMkUVSTP7Z9curJ1X4B4mijOaaVncJsRf5Cpt2KyZ3axahGu
VJCO4KeDgXKjles8RbqTj9gSflzv5NBkZm/Cm1RVf9sMw+++hQ2mBepZlh4fUblNubOoNG4srhcT
KNOPwMV/bhqpMdb5OVugUzzRwLYH8BShjLVk3hyvNWvGiXm0hnfu+3vPE3HnFqT4PQxUaglFdlcX
aUFNvzTugf9xcfmJvKjdV2bhWpwtNzgHl+qZOB5qf1r1AAlHdnVg5T2B3LjDOJY1obPaw72teddw
liN8R1bqwBALuTSPyVG1luMC/qvFQVs8mIM5K0hfESl+tPrBPWl9A9zUbx6Px7a+Gwh3dhfGcL2f
Jsmw99UKp4FWeXT01fkSyEN7Xw3wm40n16HcBfNsGlgGOC8a+ujO8Kr1HaXbk2aXAlM8IyfyEL/C
wY7T6us75myVoCSbl2rO6+UIgHFuASOY8npivVMsBgB4T7ES16SvfEdgdHovlb+wAvm3/bl7NVu9
K4eZYDxFCqeY1uTs6hLhBznXQl2PZa0UQGvwgyIfEabRBfIZOrLho1ClfU6TpBulz+JBOPMCHGuA
dHlixMQ0BnSEHXhXmEzuNO3p9Xt631gFIDZj+y/Sgw1KwZrsphL22cisjMB1971qQSUbUhavNVoU
25hQKBlBOZf2+T64tScxUMENa/9WWqDYBKgiBeXU/3wBOg/B7r4hEzyeUH736ElVFovKOifxlICP
4CJsxVtbHVKHEx8wF50EQfR5BC/EM+7DC6yQyz5lbnb5mcGna2hQTHy6/YcYhR4DuOKz8IKRaemj
R1dmen2n4jpwkffRSq21Z3HDOmvY1k5xMWQ/vximOrUYAUmcQoCfH8fDODXdXI//Oxa+++CLBz5d
tk4+6/5lun2pNjEkLZaVQjDLwSaBBCUPTr3mKGu3Jlu4y9QmhOwbt41u9oCjm6DZ1dz7yzTc1NNw
Q9tnutqtAvrFncU0/a+5jzS9+UJ2NUZzwopFOR66N8coze4vkuWMmOEnyiiaETw1eDk+wmO4ihp3
rLBm1QJzXOheLJv3U/wIQ/Hm9JUuV89HWP0KGDLLY7UE8gAz0rOKv3T6jLv0LpxtJnWQMbUsX/n+
XiIpVrpW/yT9f84Xqp4A9Zj+cfM8s3N26WorsbBROTpSC74lMyIohMovBq2nuoyKosyH4R1bJMSz
1VtMzuaOAWmwT7ztQPj45P/CqcJ01I83v9xbZGGxy26ni1u2kmHE4alGrHzQJd5onO1tVx4Crf4C
YJiyKqzZP8I2J1XfWVjIdhYJi0sOiY9OscjOLi7SWpyNaSMxEizj4sCIEnjwqaOwx0pupLhs2yM5
E9988mgTGjP+MbxwIHZ9eYyyki97+k8z5A7wLmkr42MvKLivytscVdF70T2nd4jVCC2GUt6IbfRQ
XJ9NqoXdgxLm4aM7PWWkXqPaI4itcY2SEOEyjy4vHSYNRvyrLhQrDMARxzeABvImrrKMdRlr0Wjn
tyLcG7wjKP6NulQ0ETeAvPyDHftTonXFWdJKPsj8e9YsPPyZD4NHvkrk16TCmZ1yH+bu08sG8heB
cnCS35JRl1oxJi7pGS31zW4o2+vbjlqKOIgXg+03dGelPZl2Zygfgv5V4qvSZS1F+W0qbv98W4Ad
SD7Oo6q1WgOOlvJsVHFrJIUTgLijlRHAAbTK4chV2nCbCD9vfv/8P8A6KZvxwnEMxKaRr+M60zKv
f3V+LY5yMYdJhrdJW91FgU5+EbL0L0UG5I2Um8R3ig6D8YCzY7oMZNHjR1L2q2uonyisD5wCAaGI
rqaXxFSvlMYztln4UtTWoLS0/78ZAbcsj2Vkq3+IQkd30yzpCERTuwSfjJFyJu2IA20oKUm0Cpnz
yD+RuiGVhs8hjdGIB9+/q2JWCTc2jm7eXEmFMlv1AbDovOk/b6YEblTPEplJDrEgJGSKLZU+m1km
Fv8xxC3vO27PRBKAeEKFB7D4j+51JOd/ECEJWCa5bhR1nR6BJF7W8z8vRXDytnmK6VZa+6W9ZSH3
CPMcsOWaPX08t7wf1jmz/F9PNLc1qEKv43JrwSIMBcBZqm5+JlLFUD/Nihvfn2t4Ji4QzRU7wL8h
TZyvVPkrC891E1VoBZXueBvZ+JPufOTih9pa/dUCVmhhchSf5l7o1dbMQ3BrC59HIozOecCrJfjf
TCgxKG2rEdZJH21TGf4qyuZVpVpDyK0TlT06y6jgx/84mbELkHYWnzsLvWk1S7cNCKMxSWxnPsbJ
2qSZLMeS88gHEKwlQvRie11Fu4IfZcVjuwkJZ53Zi+xhD4+aHFjlkt5f7skeGnyipG8RYCCZeQUz
ROPzHeA+k5dfkqblzWlafRZagHxIpwjHaiJ318WHaS057sISsYRrjZ6skihEeMfge9izbxx70i9A
6svG226/Fnn2tgXoU3oq8jCPfjHxxnpgTXZUudNMBcHUP05gcSaZlbUUZt8HpWy5i3G3h9pRx5Mq
quD79XbBKEjQ62mSBdfRfWi1PZknMyANtw7qRebsi+Qflq6XCOH7HistPjmgKByPh7Z4xF3LJJDQ
fVPHaF7hqkmpRnHQNhUEfJMwE7R5IQiNpoC+P7W/pd4heGWxU/c2oC00szbsh8vzGb8jXqb7AnQl
kyadH11I7lfaIcadGIIMFSnosGNbEVgcF6tfRoUJxSJkkLt+JPlNFIxAYD1KZB0Iytn0W/336iPG
mRsGkj6vsu7aHRah0S3gpdO3atq2NvDBL6B2u5ZxE8FhX0HO52IJGHlxwVli4I4EFczevNlK62Pp
c0HMf3n3zxRD3NyJlF1c+ZXpqG4hTHh9HKF/KYM7DbR6nfyEVmowzhIM3bhUW8dQXMJ34tDtbq6e
Ms85frGPPM4yIwpFVrFGizbXhC1BhFmqU6IIaxkZPnKkWhG//sDbmmBy4s2jt9J+zzxxuOCE++2p
lIp2ounwUAatoSWGIBDynivXCKyDx8PktO4VGrcaVHnb/3Ygh+tzqCg8RQY4JvoKMwO6uqE3gPnH
YnrHWPaviforFAd/XNCoA8mmhwnqMJE+3fHyCLgbAEQLltBlrp+gXcc7fCzg2cCsSkrgjo1QLhGK
tCaauPdcPIwEiEYSo60By/8zne7BXel536KpvIg99JrMgk15NFhQr5jv0uCgRA2uA8AKpSlbOuAs
zu27ShRHaVoRCAy2mAvpoI3EkVLPEweSNy/xTuMDFfxpTyGAI0e/PAqP0nrK7huPbmKtUYiXlZv2
LxanK8gGqArBaHwYGQ4dCIapaqH16nf05Ku5z8McHV0FdOZVjMm7y4Cx+GgnnUtjRjkXjM53loYa
fzgLCBvh3oeqXWybTmARjg4X9p1RKJp4UfFFD4L47vAsNMcjZT0bNv2HUyu5tCTGFmgpV4a8TkGL
7o0Q1Pc+bmLkp+alTOJKODyiZ/+3Di+/9qMsk7SFeyPw5sSonEsOXmGlCakP6HbDokgxllK2QriU
DZF1YQu+qX0F6/lvKTqkG6sh7JAIY/Wzfz8R9R6S3OuDHEN7vpcNdeCBLlCsha0g/ELX1egyLHBk
MoGaU5fatKzNIfJpdVXqmPNzUYjx+hfWsPgjuN3jEOCSwJJJB8lGpt3FHac4NPNzt29a4bD/KwJN
bG8IFzUeI/VlHBZGFboHHaetGC0ncXsWeWplhYWhXuzupsACQyBHTGnWs3vd4I7STeACOzSw1Zr0
+FQJV0tmtZb48ghiqCuzFaXxvPadv5UgcVYOKmFHpqW7hkcCy3SBvM9LZP7bsFCg1LB/blm5CF1z
WOntfqdXJ713WaY5gXbsA7bh8VbqF5zKKUF5VnPPWyDcB49uFuLtKawVm1KB9NLn82lRcF6pEcRY
huxe7C8UtrmyiK63RQFwT6/zz0hL7WVFpKvLGXCMCbc49zvETDO8KmQ6ClccGaqHd7YnGZ6qTcEc
jtEMOEVyHJhZsCXrpXlaSWstoT5srWO1ThJJ2n7Wgkynw+E/+6NmZQAMd3ac4OtEVKP2YGFmr1r9
MZoXbDkSztDH0u5ZbQfaaxFPMpdO9EsELwlAHdajN1xFsW/NZYp6K0xXvRs9iQwgBQfXnKebawKd
TMlrlKMiM2smNKjjLyU9Z5Szl5s52Kbxm3C63nWKu7CqjAk0wEU6ErtI7CuQ2LY0Fq64x0mlMOaX
psLRvzyHiPXnVcEH8aaDlc3wUaU2GQ4VRddpDdbxJoMjKOGJE8CN9ZJFFvdjZ4hK6Je35UdW8iQV
ew21qyThaF4bN3O6t8yiSkmYQ2dyHI6ysm2QFjocSdqAfh2QX+sNe565vTfBXuiHo+BNMRS6z4T6
1xxz6+I+I2eJrrcXlSCHm45Dg4p3Q6dzDO2GrSIcL9T5OVGAXdd5chRvydT3Pcx1yoPQoJVHwWib
A9S+5J1Ofn8LuyWcewMpoMLfUF8irfsRIPyDToLUb8UTc7pQ5V7U756A69ELxQ/jQfBwFcLIzBQP
5W3LKVtv9sztJd/S4nIppuue7UDwnbZ/jw+Bnj319+/j4QeVz4t3RuXFWfMJ2v+rDv9hkq8rbIJL
9fRfN30JnYvt9uAKvxucF8rGNVk+t9MWjCU9Eb81N+w/Gp4QesBaaWYiPtskdOQyzI04/l6LMXI1
xQSKwwDZndd+7g3XcF3QtrRxosLR7DVrDfCimTi1GE1xXunIPSfHCE2h353+XcW+qsd3bRWH71Wd
dV1DrPo5hrw3c41i2HLD41u7yZUE+LSuWVBlSpakgRLFZsskTc5UvqtnngiK4bCS+GTuYQ==
`protect end_protected
