`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
djm+Zk9408IL8ZoIH+Tgu1G7g+cgHmME04KTmKlBJ710HcLIFffS3EfL4C6mYbTG8KsmA2NubmvD
pkeBKjVEgQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Plp87KR5UwKisHz7hE4kX6Hkf2zdZzBJcgTvrOB0ERt/IK9vaqv5CvV9ZnHqXA5pjl5b169g+Kc8
NE+ZDrwt99fhEqCOEl3V4+zMz9DMUkuGdJcEC5gW0VSucCZrb+Xyx3DUQ7wd/JA8PJFg3niSQ30D
h9XoEd4piZeO5qkEg7M=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TvsHLTdfgVxFwv3a3ccmi67lwskNFAZqsO649VtKrOC7kGOXGAwibrtYj38Qs15qdPKCpvMwfUNO
3YSBH4kgiX7c3oxF9a/4cdgz3xcO+Tne0tkN0s20dqJwHTYy1cumv33YmUFamtPYsjXv09w2eisn
ZM3/QEH1S4qdS8hILJ5zKW4hYgTLtXze2PDiQefyF0T21JmgmEG24avziYAMgPwXRZVwH7n6aliQ
ZqOQLYOBzQIQwqmhWqVh0VIGlwVD23mbJmBxsvEsvHUjPFc+V16HXJCeyg/K8+ALhRpS2z4GfEEI
6OsSzUQEqkhUMHWR975wiAfvEAfW7I3qzqtgQg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TiDOITxRnJ2XC6rmmZ4UwX9bAeLLmoquJnxrnoHuK33neLVIgE8DyQZ15aPnvB8tYyMAOCuTBY3h
DtUQd2m48sfKaSRJTS6gIDhaK6kBpGN96W0nR0CPy7q6HE4/Q2gSokC/9ex3qLdCs+g2u5plu1PW
N2lI+paO+ey+wLJmPaA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qiA5GKwHwA0zKHmvSFod5Thqa8quduZzl7jD4ytThKt2KKIVftfb19MlkIPGrX+4ZVP1CMXFyNvR
yAp39Fr0Py4lgWL9vER5zvl6zuITilN10nSEno6Rl4NoV+ghT7Zy68+2GbfDkQPRuw1Z4IaBY0fK
k1mGCiavJlhKBpn33z/W8YzaU7JS17kDxuESy12SFLDTSgpWVU3eP6TpS95dHR14sDC6sBQeQibO
0uLpTPG+AJ+d5Xj811Gj1BiXTTMIMJS/SIfIwpVGbyosmA52y4TGQ3IFpGK7gX/vieiouK47aze6
/u67HrKRV3QGIArTpyaJfO38xgkREnuPXn5cpA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7536)
`protect data_block
TLOSykouAUhjVPYX/57wxvDv+a/MdJ41YIEmsYL1p0Z5mkalgriYWvcyN1xBgWFfV6zaZ2/eR/sx
hmgzBLzNnhKTP+4fzxhZ+yHHmcixo3on5q5Z1zCMCZED23c72mP5adkG7ODMEAmkGgZAxVXL0QMs
sKjPRbofS6XaAeTihDAEc/lXzAo4KJNAWFBX1keHPyrHqPdcBVPa9pCUknXAok+doXmvJKeVTutR
L288VTn8JjTfdvh2e8JoHuEuM+4M35S08V231FW0Ru/01ffITpZYAbVZnzI96cM8tZ6PfQ1csxXZ
K/WsfxBS+l5eBdPfpa0zX+wcnJ4dY1mB3y1//FoiWdQoPvTOzdhGJbDIOrjBLXWknN06BGPf9Byo
j1vwa+db0yWGjf1ZnUTvP6RKIhgA7WRg9ehoiyi9kdc0q445CWJqvaN4wwl/aziYioQKKO6tAfjm
xLrOFpUjiahD753WJASxflUtHWpwFGXShiYJDtRcUpNEOBuqVU21jC6oSepkFv7ONJ2tzc5xKCT9
8Is7pXs1cHNDMASh7FiPL3XKZImSzwmc4Ddka18WRr6Iwb1r5cGN26AcMevRq4dpCiOS0GynuiPo
ILaK2xgPd8IuKbmeT6KaTujIomcTMg29irM8ObQd9QH85h+LKYssBwPcbsSuU1u+BYBxHKEQO6nK
TdxSLnAq9fvYRwnu10Aalr6Y4qPpgtzV17x7FbHl7rqGs2cBq3lerSOOcAoRbJA3IpAkLGzhzc4h
E79LFc10Qllqz58nd85tYUi3wHiBlyAn50GHJFUjtl+PmiSlJo7cH+K5n031baErI3zLCqipl4UL
phcNmENVSdt/8HBbsKk7wyd8/Kup8smpC5KuWhz+yxRjh9wX3uUNjWlKy3RwXeS6p/iWetzii6NJ
C0lrVSpyoJYfFDRohVpRVrZoFXxGPM6zCdsc4IChp1Jsm1Ntm+Hq3p016qzURMeWYRyZlkoDxSto
nYbZ0EPrPmMOP6Jdq7+9R9baonVEhKtNPz1OpsqoOlo+cRpCdA1qAezIWtRLAZGAqswjXbQm2NYD
UtwGpOUTllCdUCTjhHN4NdsEhc2QWZQN18XUhHwNuFoQsIGu+LuXIQMbVUBQ9MK7zomi/L21Q7YE
JTqu5DoRqwn9oblcFxD4EkYJlklacrKzvendmOJMWIeuwCsyOM+t06YfWtDnms0vD3x3xsDDFxEu
+Hl+niyVvigoy3AwIA6Qs3E0U9X4Tl06UxuCSLmsCPhfVGvEAXvn6Y6y/3BdVqmYcPLMCGUhfcWn
FzoH5S+ZWj5PJVGmVnnS65G3sblj60XiR6NK7tEjQJKPPFNFWOzzvK3VgtOmzQ2RNN3cWZ0SIwRT
l1IEt8J+9njpPbnjD50OHe5/YD2P90h0qKHrPDkoy7wcjDD6vMpbztbduju34ywfMYE/kMQ4ZvQW
MuyE73I/MPJ0kPSk3V7yiJv1MP5q2lDpwMaI0ll9Lf6e1eXcXvs+eTAPSZ7qO1yz5K836DaeGjaq
D9W0hp0PWwg6NVimlzyfS/Q2Oz8C0W+zwNhfCrUAyGAXHiufu7AdbPUqNT5asDhanKDsztCJa4fB
UQV6Rw1NinvQyvYmDMshXILCAp2caO2pItzbhgLL08ZZTjPfGOWNP1enwDRDrinx41yE8H+yFdi2
H0baMBW1d+DFjYAuzl47U0rVYziStUJMKnxZ46mnajmf5e2j9l11cNCxhFeX5VsIFHqo5ca1C/2i
/72nZ4F5peIshtF7fgNbr5yAZ5vmRyXgAB2NrOyJQGtbRv5jP5zDtsR2xVpfXfvvTPBgAZawXTNd
YPmKCCGSYgsqwholI/vb9MkfazT4lGTzVdYSZ/jj7/kQ2oNh7VDk3EPy0iCzDO9sSaFa51fPcJNZ
4HM+5B/tFezR7RR0HR3J3XXezdc2UE4yJBC3TIcBW7gEOrlnPhkdWKkAqTSm0+b+nrseqY0ijxcA
Qz0MSJ5BHlhqkRXeEjvyuwQJr95nOEmw9ueVRGzSuO8wyZCEeoUQiqm80ujOKnoaP4kqun7O7pU/
HEP1c4AUq/ou2X1/nJCZ7YEQFSWkJEdXVRQ1VVGZtqjxnJspOVzjM+slrmxIOncVvRrzyFeaYCfE
438ymyB2a84Yw59LhzW2WgsVofua/B45CYJMGL6+BCcq17PDBlZ0LxlIu2cUW6glPAXENYDGcT0C
6ofW/z7ZUhqS6KFzY7v7N6oRpRG3FMngDFBjwbXfL3mtPICUXwSdj3h/QuEFE7jAFR+u61VvBm9u
W0KSX1Kqf4AqT8kNnb03T0ZTo8TSN+zMAxl+QlPRBQwCatU2sM+DbqrOyH1KlRQubp4QhMcSrukz
Ye734jt4F0ZQr75Mlq7S5YaTNv/7l/jve9qjV97gWe+VWmICOTa1SxM1AV7DTgaNtRWpRLBOQ209
kKeu1fm4QvCuKG3JBEukGtWrpAron349WU+LgVGMNxrei7fu5qAl5ogXc8lgHpdWXG4aDQKRSx8N
V3Nb/XS8fWfmNLL/vGITDmnD07CcQuHHuZ8gFiGpuPJFUhY1nmjiqDsAauBmRSLqI8xd8Ie0kuVJ
dz4rw2dKzy/ay0tsv87J/fUDcTgrCeWhd38WLocNvCWw2VaurMPTmlM4lyVh1Mo0Om2XY2GzJYMy
PzEpxoqv0lefoV8wPnaPPdC1NcUyjMqycJ3TvoF517OoziBp6FCUlYkllu+MBqgmXu9QoTMZABMc
8i0AS8O4RiAcGFWhV1INakIr6A9mZjs6AT3j2v3CHGFRrtj5l2a/iLJfOgjwnpzu/6Ndddh6RnQN
bTt1bhnH27Chc/xuVx5NR7ml6nh+FCFwK9xNkyPaCU53udwaSK+J4X6Qw44vrWw8/rqyPw2bKyD/
36AbNSRDHBUMm6cfqlRIOXvxzVEAppuFD4uwuY2BEkZ3McJEYTdPrirOIhvUo2tSnbJVE7rYx8yj
EYdbyRZEtF4G02w62/Aa+SvBODfjkOuHpXHLsZ5QdFPVodF+rM/shIzkHjhZmOJgJdGvrtbYDWd8
alP9UgZ+jwm1UyWRVcpRK5yqOJ+0FOWD5prnaq0VQ+ePUGJ+B5jkqP68l6PdmOo84E2DVvW84SsM
d5V2E9aeXTZMXBI/e8U+J24TUgp6JyGeUrU60zxc8jZ2cPicPpm4XEKq7yHXMoxHmg/movVxBobm
ycFcoG7CifTN84lqccoTIbVKuBWRmBbCq7LFlgpVRnsQbxpy47KDqHCDBm6tfPuXN3oqJXKZsqbb
F8YnDTnt32uu6Zt/uP3nyjEHGh+B6AnG/ryNwxNi+JgvmhguOHZVnx3sK0dhdZfU1mFqGAv6G1Cu
anzQMbwHch6gXf2KihT5ObI87O6Cp0IB1DSfyhMSxg/KI+cSBI1BgyoSv4bBpk5ZGoPP64lrXw5q
ZOSjcv09qcwNxkKEbOWxaotTSZKVhGFEdxP36kuZT0GpUDPKdc+Xw5XfB7pzriICqt1LXkWU9TeY
dwQDRN9dHvUAgaO0t/hQFnXBqZN7rFTvZmUwqLkRjgXmEJw2NZ6u2CUowkUZm97FEOB54zIbNgGz
eZ6BdBxV5lgimsdo/AfL4yZDtCr/bMTkEivVyX60Uze4kKrUWGqEkhFcmYJnk2uzBZjyguLHRTbn
syMRpUER4zXLnDCglV1SVN1Nqn5jbHvVinhgaPtXLGkSjn0okdiNjZ1kkk0gR5f1GfN/2he1NKCv
mLdAQMfMHjIPTg4W6ZSCNV0PcxmNrBY/uoqai8jfM9KKRtOciexVOEEOiYUd1I5eMhRpnnwvuKTf
xGtSYqWtRxy8JCxY0Vc1l5MFjqtc2Rj4Poh4PVbj94GdG7GcnX5r9l3pUnoa6Lts6qQQ3kVbs0Cc
mKFA86tw/KJhLJoPBEL70+d6N573iNSomZGRKdVNKBsF/ZGFZXC2letJA4PMGhxz0EHwTyRHVBIY
2X6+zfd/dcnjtTG34/qMPy81zqfOmsjoSa3JrdIB6QYR7C4EsQPKBhGAiRHlfHo/RGo5f71G5TVc
+pKtIqwUpoPtH9yqefCGoFyTUD5eFmX0r/YmA/YaFxTbtmrIi+IlEWn9wUgk56LugPWhiEA0g6BC
qK4e9Ml7mi2NtrIG+wtsYXsk6uFysTKG48ZoIwJPxe9AguPVBarUC8RUW2zpqSkYdghK7QdLmL+H
fq/sODb1IorRfN/cpkmp28oAR0beRLQZxwvbYS/sAk5eYVYIN7X8oc5hK0KMNnVqxCkwPydSpVAJ
Y34cBj8RVQB7tLm+mwiDwDLRQ+YgsgD0Nm6tcddIXOBurR3jW1AaBPAm1mR0qx9LTDIGcMQhwaa7
nFdubCQ53n/UDdW+7TAR79we5IK4A0DL4fOIYlVop2oj/ZZox6FVo8c6aduOKl9QBZfcTV8kGf4b
AyYMlSJPaX4SIitqSuzeuzZVxw1LEphXhndaun5mlyipqoG0C9s77LeAdG3+6ce1lER+lqTD3gW4
Y5xVuHxQTF+Q6PdPobF5qz5PAO7sfs6vkLbDkNVVRqTG6O9cP7pXjRhWlc2D9PrKICxOzhQA2yCs
Q2g78D5DQ1MPj580aKeqkmhgsKwDZYMMC557ofC5qyYg+s0eu+FohX+Ys6RHW0zACYfosbnbn8HV
5S1va/0ZrhuwYsagXJ6EEU0egbCo7PPkibBjT3cxp43ewsVHCplKVmUkdXs4DJLV4KgMTffnm/PJ
pgQ/ceKe5QRoBw0z2ck0EB1y4nbvGRFffUHDr3DJw1JAfCA3pmAGxcCWo3sgQss1UINXCeqjTvOS
ZJDPDpPg0mJn8zUkW3loBzWvqKeJu9TD58JynuTCuO7+kw9Gt1rUBrBzKuSB6SsSQcdp8qVsaC+q
Ko7xrXdKYDgs/GmzKlcE9/mBOo08r/NOiMKc0ZHLf995yJ1Iooa52p7knDE63QW7L/MqKC9Uokfu
NajJnKPoRbw35Bg7hlz+Ji5+eM+9O5Nt7FgO1jFPoobZMES8gPArOlI9BWpwl80eEGg73TrcBMJi
LxnDG/QpJDGrM69ROGmMmhADgyidcw8JMINNc+YAtV0bOorw3W1UWlokk920j9QHeWMTM+uZ0Dal
rZUEvaWLPGw9Nl5Kv3OJMKHob+vcFuyPd0Pa4W24em7wGZwMfJFrB8DxhGiX5qk7xsmc86OUQqur
caSYySOLnQgJ1oC3IoSNaCKrqYFMkKu8fE97i2y+hZvRACB8hxH3gsbiihhHoxpkQt/+h0m1ETbG
tN+/y7Ocmp6jq/spiHtcHCobwGXnG0Jemnl5XNJc9GyOeDPjhqQYO3DWiiQQL7IhHtXSU7qfJ/hm
UNZvB2qc/mbLKFIBiqNvaWBwmXrfDEM5bWKv1LRfbWBVSOf25UUGDwGl9XO81QxopvEJ6dSF5dgb
7ljTVbkfJkh7zvyHOFkc1Wx7MWJMR7ezCgVelOdmKVnGpsTU/cfJI6u7iR7VJ7EVtx3iFi5ADQWs
y+yg49x8xcYVJ5QH6eJbuNX0leT/ijZWtELsA+C/X3UBDkWzZ6K9CVkLo5ijld42KXsTWrUFU3Br
KsjcmW9dwNDozzTey1uENJP9SxqHk0aCvQRm1sf4G/a1pDec25nlAgeva3KUeiOE6k6ssnzUBBt9
HWclLlZ0jGUvgEtpMuu5TMk3GoqfGLo4GtimJVbaQum7E9hUw4agPiPQR/I6jqA7bKZEEAHEVNCo
mDorYjLvSG7pcFOWGBZ8zRJqMoxIuxCA0UxkXB9G8hsvRb9PMAiKP/KIkxtm43xwO1osoIGx7ESN
dAyoL0sBCK+Y+1Wzc8QmH1LaNNOnmV2GJsWJqmA3H5USKBVB8lJoOx2/9DWncXcqdeTxJbKDgcXN
k5X45pe30k0Gc3EjjWNYjr8ZCdsrJgg+NUMWICgIEpash/1tP5rUdit1Ps63FN045kHmEX+2byuZ
zIPbn8pwDgLNh4dj+TcNVBXsABT8DcFp1bK5AFM8MX51i9xm7h7c4mYgnt9zdDQBqlRAmGRyruqZ
kIKve0G6IZV7GN6sic8i1cVOXVHwiSu1YJJAxHYpe0OVWjshztApbN+XelI9qjCmSQEdbkvQ/Wrg
8WAzGfaJ847j0Cl+fpYvSVh84Do8uZ15NeMTGI+zHJ8cjzuz/4HHVZsbCd5R9/baZM/jHIOE67wM
JwrmvVejQaanpFsb2/Cm0NCDtOCUQZmLxenPh4yTsRDDizHd8RIrplnDHUpyi0fmbh/meLXHBTic
ECohgBiY5IcBhBN4bQTYsc1Papuo340t3MicM4Xyk+MOg9vo10qex/+ibnlEzUVQMiaB6oCN7oQ6
aZHa56ZmNZ/hFs88LYimKg7RcFsqeD4EQxb55n0pStNVzvSxyuSpcjJlrAZXdp8TZedKJFzZoNyL
+oYx3zDRsVhP5gjhbbqfKgoSnwdVIMKVJxa3EZpjLcRfWHAToLJHIVjDyTS4PggZS/Rb8N4jHMHc
FUSjQg/SPFK7SKLZko8T92oFGX85+oR1AXZBVc93XaufHpKxahdIBa6GHa7VgZXnK16R9pI1pYY1
g12ChQOE3cUNINKteHLy34y+91cfV3Ih+2zMmxfdQf/Q9lQeK/maUkO01iQam8oo1vZZBPCOyqfz
ChysP1xhExNYp1PWBwtRRmmuoSdbg06R0ZJLoiJHodRok/xRFTRGO4SdgiBAyzMMOUnxuIwWxXKQ
aOu0slN0Cjhhb/jzsr6CIziXwktmGpKHdMbUsKo1kHPF8KFfbLyEW+a3qAQgI2rGjY7EW8QI1i+A
3NbFbDaDKLKAxkjFqVhaCtD4coa43Y7ahf20tiiTEyp4EoxVYZBx1pluOCC7vC15TWWePAQ1WNNf
hy4+PRMdFOSbmC9QpF1R8rLC9aYR6zFXXljxoOj2NAJZmOuU0KTXycrYvSeQhfkM778JN9n7dour
oIicJN+R0e3I6tqXJrYjppUi+xct77c+66wAh9pD2xficHq6N+sWcUqqV7jn5XPLu80lh/ezvojM
wKHmVrgKzdHdBS47PZ5og4VA+OtwwMFJzQ3JH2SamF9mHIP8ZoB+uJ+sNWm29mGuQegQApDYFajO
ql1aVrN3B9mutf5Spa5bDbx3/RDR4h9IRm7zyam9x9AGqqTy7rAeOC7HGhC1W+nzrS3sj9zMHCLS
7oCHKNSnTn7kHaCbZKN5QLkin3Nvya/YWmdHrJiYWssesYlvYOjq4oydCmB94QUx+SVz0MNW6/2j
dQhlAU/OSmMWN8VWR5BozfX5lCpOn24HH6QlTBoqQyJuN1dMffb7yeY58QDPnDNmNCbryR4mYYuq
Xp/0bLuRWK3+U8te6cR5Fw/72F6cbayhXn1WPv/XwGyoazp3pRLSeNA0klD1z9MGKWKQKCgrCuOY
WrqN7Arv3RtcXTPvlssIa/eRnJT9aZiZgOcTUREmPA1e+c8xIdLUOZ3aRdq9/kv9NilZyIscx5Q1
akvwODDLs6OiZCpnWRAxP8PznHA4sf/kg7QfrgkJ0MDKNvWR66JUJwfo8YPCgvR02a4t/NQhxzH8
RGzlrje9a0vRlq4yZwDfGd5T88ksEkQ6ThnI4u8m8oEgmGzJ3IDNVyn6n4QHjUC73tEVy3wjQtbB
yXCpYWXdNKNdqkmKvSjULyvgTlxmTZDt3boCemP+JpHEgvFjgz5N0s48bRlLpKBt8wdpHs11xwE+
jq+qeHL0vqYndOSYO2aYO3n+7LNOR6qY2d8nmRk2n8QBdHn8aNWeRvNxSbIgjGVhpr5LOm1dp/Rh
TqPGaGYa9Kzb4ttnQzfKKrMTCZfv/2sGZQCGcfm3GUvPQRCI3LUWx4U5vs4lBO9ABDXBPNgY5ZLJ
tfDRms7eu9ZYN7m2Wgc5YNxU0OzkAkBdyXECvrgur96Cou9vtX9WNtNZ+GN/lejK3rkUg/dwtRkQ
xEBN3xrPHkw/DHk5TBE0iRdap1SDgR5027GTLFUvmevKmerTHp5Y2uoIxdhxGmMnYbCSra9HjLuq
LW765oFo7TzN3R3m+teIITiSgWIS6Xb1bH8Sm89QA2gVsSmAxEKQwsk2Nuywg31mjdHnLolk2b3r
gL6r6YqsEnnb74aeURvNZAQSBNK/xTlUpKZquqXi5J8+BloHpxryvFz+K66ZioAs4EiFI2/ymQoe
7pT6s46gpIJPJe2GCvK7hGVDjTqUHoRmdIRq6MMWjoxEFXSCYd5NfWpuHastoq7PUYUznC/9WxQJ
WzRkOSMp/XLM/33NZXBMlwuHwTBiQatM17BPcjCeuanq91a6yj3ZqYHvanJ4OzFREBnWGtmU1XAm
8f8Ga4VqoI39BrqNNgXoqBQVFSeMVbQsqjVcV8IuVO3tRmW1j+4xO6/MScVPqvoapjUMvpJyMqxo
vZpJguP9TVwPGnI2F4XecxWWvvwWXrXXf/+FiTaS/mol27dHp9e/14DrBjnoOZ/bNH1Quqv1GYRV
wJSHyCNJS3Y1wZF8QYspAi3ULuOLihi7fpC+TYQUQDMeW3akcDCgCra8KCoDpsgqWFA7BsavmP42
hYZGKDLCjwcmkPOeylwyhCl1PASnAhQcfZZ6s5BkkTrE+pm+5Htlz1whzE13XQkxvtWdhsYp2Umb
dprrxD67DH6vL3EHJXAwK76WXomi456wKkhcMgTSZMkQVQFWTcWqNVZqwp7t5O4O7C6nNZIa7wg8
1jGYPpy7Ng+nV8DXS4AG0SEWTvIwfGxd1QEuoregrG0IYF+D1hu4kif1eGDaeKV/qazJimbi3p+i
VmGJy87o9yxF8KBta7j/hKFAP2PYLl8e3scYNDX1Vdr6xVSYcOzDiJ9pj9WTPUvzFdIM4xPNe+gb
ZVAA04nHvHeGxrZJan7X4F2dPIVBYYaQBPUK0qLPafLTay/Rn3e7RLaTQAo0h+EJJP0FqADBsipo
TVRmnXC4nIqkUp/6U6bOYIMIDQ6vtA+zDW7r5DmVpZDJxnKoYrUCjgYEYYkwcN9/PstWodjvGGnU
BC4LRjQgb5FG+0cis1SBT0MyW7XxPBw0OItIPoKKepLfqD1IHJrx/R154uW8FHI26Rk22pohvyhA
hvDTrKKMJG5unBrOU+Hac9anrl0zfeA86QcWR6OmOuaYWv4yp7l9N9m02hbkRO2SPudO0G0dD10V
sCXm7fT63lkbQrIbKEAitiA1Z7fUHZZcS2PFxkEg/zprWw6dnqPiKBevbyF1bfDo4XtqH3K43KJZ
DkSzABQFSfNxxwkB869VqQy2tc+OaUWurXjPvUBg8rvoolSbBVcwdS2f8CUG+cXvrGozinpz9Y9G
AHLAUyQ9LvR0u8SXtrcm2ke8Pcr76/93X8W+3fsBQEfWviQyAkXk1Dky+hY1wUvVRWt45sO9FLnc
ua3+UnqQjP7RHHeywFgtqAW/SEHkV1ydPAR3xdKlmtYg2Qez3n6QTNq/JV2dfnTBpVpxopfX/o9q
PeEhlcefrpuySJx8TUwfXME9b3hrQYRvzLei+3NUnpRQ7cENFimgOfhRcWCgjgnzgBYmACDJCbXW
E/vLCT2OomgSbv+tBDqPR3f2s/FyqsmfiThMcRND/4gJIGXieh/tvW9dyZqGAJFcHwroKuPCLsxd
cqSnKdjSxX68kOWi4ivs0naic+C3GHTQ/lsXKJ+lcqzt+YXmugGDSZYJE5CakostCnFc/TvqWbsI
Ilhz3ODGtHcA18icGyiypK1NBpkscFSSySl99u4xjfnFkhw2ORBK5o30avp677aWEXAJSj6AsRrr
QP/I1Rswm0dX/AHgiaDAkFe25zRnljFP034v4ZTJrb5GupZwXZ3IK1YjC/1khsFp4Rm7uLwBMlK/
H4x2E3G867ef+44ZEYVEPzELYW+4a7KlxwRhtMdKS4O0IGLL0Pu5F+KEZ/mmYnPhcksmRmjsBWsp
+9H4oC5KHto7TVYPZv90fUPo2w7vROYTYNNpC4NLBCsCdAIKnXGFuyCZ4k9KkldXH8hYmbmlrxi+
tixwTa64DbHa4H0xZsclrCJUbuwkmMP6RHN53yvaQhe3xCXVAibHa/sHxQbdrJRYEZhbN/zzgFGA
fiebWIMkF7bPH5T1
`protect end_protected
