`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LQescFkx27XclDaXvRmW0O+G+YGbtckM3Txzw9YSzpE4En9K6VeB0in6RayHDk5IS0l1qsFCsHIn
1kQ0issnTA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fez8qkDySM8AgcB1U6Pd12i0f8Pd6yPtqxf3wVVmyd13quRv4gyAlXC/jnf1tJILfsk6jCuWrKCY
HPdeF0Dq2FJ+oQ2Y/74w9ujCf76pQqXqB96f3r7DJrDrCggxS0Xn6197l4quqp6wcvTZix86iUEv
Z3iYfLkjdA7aCNhDVeY=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DvJmj5x2lPPKpbqDEI8TiihWxWOdcT5scUxipsJ0GusEsvul9bdcD6lMtpcoAqir89DOmCQ8cx1F
WJUIfd7o1ncHb8btx0zxnZu3/OkrAu3xbEUbblTtDaDspO6DX9OCmtQS7EnREFGSPYajfN65ad/R
6GIQqqJHZATadQ2lcInn9YcVCXNO1el/eq15QrYeBlVown0VQtbe2VwjohUwSMmZYXkSNToc+q27
pksML6wG05tVkDHiCLDTsZ2lkIy0fI8CjEUzPMOomUezr8cfukvgLx1hVlocgw+8VGlLyeKdlgkr
VaFUFdHpGDt6fqP+bNIqAkctjrlX2huf4ww+xw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ISTjs/q2ObrnnUGvt6rx5qrXdOe2YtDoNRNOauUF/K5tWo02EqVlrawemfPne+2xQBEi+AuD91by
lbtz9IjiRsEbnshQMy8AZuLz6KoODdWeIHfSfO2T5mVMpJkOFdnnoJCZXW4Wnc6yrKGMH2EIhyCk
csGZQN/kLJWFZiAsdhg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
loMGx3v6ScmoyTigehIS52dUe2Gotau12+5VXd5I6Qw6hN6tauDP/mt4UoSXh2IVcERrBOFFOEzp
0Gfv5v4w/oewkMT2myuFN8zCELxY3j4PpVcUJzUXufMvotZg+uPQ1ZCZDlLKIzIJaW5Ou09WLJbP
eOGWH/b8bBq4PgklMIL0F8dzNt1L71hWLHcKb4o0cH8Dqqesl9F9f8hVBwLeVoEDPGid2dBdrEvW
fkZ11yweSUFd7NbZwFfJqlAY50ze6+IN6KsIhMEIcVgJkVnZhJVus+0Ig56zlUUzieeJcVAA6pWf
XQ0CJFP6VhU+ZISyVPGqmBli/4R9LA8IybVhCw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10784)
`protect data_block
Wi9xkj7CS+Du4K7/qi/Xl4+AIymkhJ7N2PPaimakAj0IPMZrcFS9Iqu+xCccR6FpOnIXtkSqSYd7
eIhlBg0qm+IxCmkYk6ezMScD5OVuoNxX2oxlikCe9XCqC94w3fpoIf3LbxIFluovi+hmyCVcIz9M
rkmK1oZP6vbEgvRuq6ILJOdO/AA6c3WjqV25fZFftvNddnf08FFeXKA0kvKapmqujrO8chb8CHra
RuSWcfugjspYbe43gIdr8aGcoPuBKIl4WXM90xoSQ4xUd900vwauY/ApnTU/P96ecHCkd8rg/h9w
KxzJ0063w9FonWYRaTgey1Y/C5pFse8/NA80kcopCjf4uhj4hAVBIOeBtMxiIkhRArxkd/cahYqq
NDV9JA//hFawsnfAcdpp/iitiQ88Zui3CkNRWIdiVpNh3p9SnSfNK0jjnG7ZPZCf61QcHNKnc7uK
UV9xvDvkvdbA91+8aMHnJypcTTkpL+hf8yzYun5JvayjkKBWQXHCuZFq+9AYcWXbBUJGMlEQ6xdU
qST+lcNOHwZjiPVMUYIGiN6LhckwhrEn37TAWQJ1vPW02dthV0o+jdgqOQv1PHWiVyapJB+O6iln
P0G6zOivJw9y0rIssOqC6LClLx2eU61LqCiXBl+XuVEz0e0JM3MGef8NfI57b8Z+doSrApMUvoDC
0hs/OKDenrDk7p/+wcKJ/uLWoiE23nioVyokM9gfb/3M+b3dHEJoq7rk5dAfd96TwJEz66zpCX0/
SuxJ8FyDVIHKNeY0OclJsxhb/0RvonqixecVcPNDxR1ChOrdR5bBbqpYBb1A9RknWxt3fjOMVWcP
fKaPZYOzsRpArPopDcvR0uft48NwBIPbnncp2GgshC62RCyHjH5U4d1SHEQ1weeVg3UWPCfUmR0x
n2zZ8TJEWxTyTW9b4KCCOCtYOfUu1FZISUz9Hb3oWLOhf+5Ex6awRiGL51fv3pC82bOLFB0R758s
IYCbbNQzHRNmpuvQrtdy29pannr4GEGpUFpSJ9oKOdJB7kJdYJXr5opjnxVrEXlwi0r+9YqJ7jtd
+3zh56MMlYGEJeswBnRT1Rs55CtDCu8WZz1aT5lD9k0kwQktTY/7/ePrr9bHfZT5DBRr+b07Ji9l
9RAjsjA4ji5IV895smf7Rp1wt5ZVPGC0GwI/Bb+A/6sL+8al/9Kn9dkwURV6wMTcbgRY1Dlw7Xu4
cT999+hXm+HBQAhgnMj4zbiz+/LWCpGRFDNVomFOaVbLZ9kM0v/OcenGhxecvlT/teDhgJQYXeCL
PSPq8WxwVLnppMomn/7nzFlviJHB9M9ei2+YFe1mZdxyFDc7Mt9aJI6K5CYUFLHsdEJ8dNkOJq33
oBr+En+/Ky1O/qEvFKMmxddZhgWmNC+zI3nEuIdk4AcfttPdznoD+mIdgKC2UzCfdhoX6xaCFoWE
kNh8glg2Q+srDuJMOLtnA7Iy4l2bsGNlZRgN79QBvEJ3mju8DWLrRoEGnndgYy3HCP+QrmNjdNet
c3qhxmt1pEX7sOT+o7MTSxpicSkgZAzuWqH+LHmNM8lmL7kT81INVKbEFGstBL0gr9iBZ8DcqiCA
RyjBilaG5bwPv2x05LKEwyXF4Vw6GIbkewO27Wdj0d9m+wdEAhK5nXI5mxY1SKa1Xw+tN4Ca3pJ7
FPWPlELrc4GkhgzCqOyijpk9/py/oUEVDPjnj5eR/c+ptLHZl+U2Ym38iX5fYtvEzhlaBpN04NXA
Mn3pIMF4daJBpBO3zqx3sTt8Efqp4NJH2ihhT35TSKhgLxq+5+xWR3PlpRqH798YEXcqJOdHfILb
VUOH2KN4ByPZ+T+w7NarMfWevux0cOOSkrWCXjngkrfkayC6huUF/SZ7Fjt2leI3E5kWypOQx0QD
rvMfu6VJ+h7E3ddiB+G0ny76HbpKu8GSS9y14tbWuDfIC0vtEMHTWtYp1ih9n2ejM85Q2zY+zLWO
g85po8nhaN0HZzRcQYviLrW56hrV0BCIQt8P8VMWl6XqORSIQjYxv52TQgK8ItCthk9mvDdAi+Mh
91CyfdL48zW5trMxiHG/r8Lx3m5iXmFDRIz9lFsoaHDibYFcV4WDBdfuY9oxc2L0q/OtLLfQdvTT
ipuKc7hqsM2y6gsWevv1y0Hv4c+GkwUP5Pw3fj7dvEcxdD5ob4kcV6QpsporvW5NUl9+em5j0PLG
C7nNgo7l+5qDha/mTublOu1m/SkSaxGfGT9HsS2hh65FSDUxU7orLy+n9T3TaiigeK1/Mem2mK6v
fiJnG8DJ/EIhJz5fAjTjy9LSbScc93QrZ7mBwshHOcgjQAIaOG44FVhfi2FNAomXIrnFYSIH62FA
gWffWn1XKPzVOQJa6txcyhHgsi9aFs092UhqkgCAEGCptKta6lzipsWTG3Belhdlm3Y68jSxZmNs
qF0nya2CvKNlL9d8r9X4r/OntIeTUKHk0er9BdEVvdPqqgtQx2d7j9xkeJ7KbtyMzHvCGxBQpK6y
SWQ3QPdXCiTet7+FHYRFcIKULwiYPbV3Xop5iNSG4j1zL/jwgGnKTH4g1Shv5sqzS4FgBhZIhgeJ
ox/iLg2cYl0RUkSMJsJ+qM7BH47viO9yc4Cx8/k1EEHGUVPHVDH9sLZsNMGOvqSii9BM+WTM6W8k
dm6tP2VWUZePONN3fZ76WfAYV3xmnznXVuIsMay8Hr67UcX0cThfZujG39QiPZJtFMw/zT5RvBB8
30tdOBG7ojLwLm3kI7Z6H3jwkvadDlVNO+0RyrxDBmMuOoQkbMEtUDVelwcZI/+itD27G6+IOOao
prObBnTR9N+Yn+chTkS1fnrqK8s4gHCwbTPeIFgpSBYtJ83OBTZsCF7Adm+h96YBDWKheAhJT37Y
by7dFoqCk2nl8NoLGGeiUEJOh4DhW2Y4qFPQO4igE19VZziuSzYwWFBmosANQBgpU+QGlLz5lBSe
1p3/ff2uB4JQwisFB+GbwoY0pqk82Y57SdhAywpMPYc4GjADDBWRKCLWQuWWLgj0AAIHN9r/nu5B
MXK5mftrI8ArlbUGdyjbbd+7AEECD5TuDUKyeu7zlJ1AgtYTfrUDuxHuYye6yLVURFF66HbznP3w
bm1sZuca8XwQpIz6wo6VKUHoZU0yVml8iSZvkJp1ke/c2bHTr8VK5KbkGSdIOZ9n3rawWAfL0rjo
Ru6YKbQEhLepN68Jc2HuJsL47qb23niNEwYZu6Ef+Cfa3btiQb6EDaxzae8d3/SERTJm7Pe8Q4kH
Sp1twxjOBOkR7rxQrSTd04gOVtiqIn29TBOZ4MGFduvHIxFIHHpaFyQE6YZ+fqkegtZG/0ZEdJom
Iu0Lcz8vE2CvY3okyp45FdIKidfb/Xkdb8qmJWrA7YwqKD6Gh40Vt7kuNGW43+9lkjFwaqgCSWAJ
7DyTOrckwcmz95iIGXFrVwhydpVZm2carFJdApfUCHY0VP+agCcmB/9Tr/UeDoJ8oYqh3s3VyLKW
VnDUPNQy/JH+SQDlsahevfk646raUZoFJpFoOtkqJ7kN2UI/QrBU1QUGIOvWUgO4NHj/iXsq6ZOI
kIOFGEIEvaWnV1psCwoDg3GN+1zj/26x++xzYqvSwuxG/tLPPH+nGbXA9DoVeqwb2jfGF4TuWVya
fpDSuxX4kFa/VrM0Ywox3HCpow27GX0CBTyKj9eL4ODWuSriBqwbZZsJnd2T318dpvJ8cgw+Zagk
p8tVRFiy5mWKejuTNKS3dcvbMhN3sdKB6ummFtAsRdeSlqpo435kpW5qemzYF9tf1MM1Zq5wXv9r
XT0PksWyDskujdNxo6W6rhRgiMbTHzYfqaGYGEb/J6mqPH/Utjao7s7a+gHSlEG1RqSzXuMmv3/0
zmGToCmozC3hdKVWGODJGaugNwhe6b5AeU4cX6H+OHcr1ZMJrb5cFU/0VK1jGJ/XhkVz2uIrZVdT
3tM8GPOfbGjS/um0RULVaZlmVh1dRG+4t7VSXebNZuQ0d5udziMvsAvJWjI3zA5UwuxbJ6ASWbde
dITXmX9QVUlu57rm/dh/ynLusds623Ig8memLMn/YafYL6obieDHDhOiclEMfLxuCVt+ZxYGpaek
A1Vwf3FC5NGkaEeQgvKkX4x029UwaYdJkqNir8PxUQl4Xc6EQcvPsFWrx1pqxUva4C1+B1ccjfnI
sPc63p5KW6lJ3AQGC/i4bW4JD3c4/zmAPFqEcd89niop3in0KZYflNTEIntYWZP7cj3xJ5Y1kY7N
D+h59G0rHI1RN9TgyPsmYQiHUhRP5v6ztvVJqe14BYvrjkcQ5nIIGyTSsQPMUVGI2qRB9WEi3Q2Y
mtC0SpVqd8YAjhnfgrD05YI9C640yq6+cMPgr6JmDYob3AXd6piqlMZMvPnL4farzStR17DxFE7Q
GSFm52YtcCu50baJ8dg76af603SrzgnZTlzOqxlHAIr+2LwLrAcG6magVZnZhDBYDlNIKZ4vfT/E
9+2sguE2BzOqf7FGy7ATB6vrfeFYrAmMubA18yIs3ltA6ZpPLgE0PMW4VWK/D633doiRr6LXM5eT
8OLcTOZsr0I07WFc4j0ST0mZOYdwSy7qhCnVaatHEcSbDivk8iIg9EhEr/j00T99vZ2egI3YCeSd
ePc9zSSvWvIx86SqotLKGmImdp9fLriRPkNgZxVCOzyFiJRRbqTwy3QiMaikB946CqColEfTnaHC
I+sB7T52TjM7oh/W+G964Nyxu84bXymFHVcq83kiAh4Tpxe+/qr+k2dYW6hJ8oQdWzOKgdnqk12O
BQRAtp7+LSl6B+Zguysx5xCBFfykLqu0wCC9rrC+FfajIB17cZmDcnLdCFgGNkdYhkAUUMs4sc72
7+7nyP80H8mMRmzl0Ge7co39KoWJ1YXzOqoPreBoby8oogTS340Is+Q2inlFBTHgQNf5F4kLlK+5
cRzVDYxb4xeT5yaQPay6EAknIXxRvLsvo9UCmPQHRhGaeSmL5A1BHqykihar/artu7MDkqBfYZdV
ScjC5XXN+sSC0RKY5hazEGIFJRNsLbwYvhZOhVxny7eXXwqEXRGTWPwnTY7f2skc+aVTl8j3DvS+
I0zSaye0d07xhqQp+/AOS5MgEulY/LhGrNk+Hn8SWG8M43KZRxL5LM+N/FtNUmMMIGM9S24n5SEj
KV2UTtarU/zJIjE5GhT3X9TdCmu+0R/daf9cMRebnJ8hW+u5B0OXXyk30TXmhyWVanVXOf3kRjk6
a7AaHiQb4BZ+bl3Z8mTn/LKOM3HMOxDV1x8EV66+JorJbRssO63vKP1h3SeR96r71NK8ZZDGHs9D
qlZUpgHOPXFSKPXcBDnEir2ojhEg7MBS3ULNK8nMliKZTbSFnckoFGDfYR41ztpDztbNYi0DDzH6
v0vR0f+r4o4jvfnrmPEnvAeL7Udxk0rx+bXF5unjNl01Tv/pBQ7T/Fm0OJwpCdWCVMPoxKzAzzCv
Ch8lhj7MEfsgWVoxa3OhWk+Vy8MPSg5sqBVB1lg0SxZAuOetQMpALJA/WNAEf9p9q0BHSZg1FDzD
PhSoFtFFGk/XX69sidpjYZFTz86+2vVYCoCgsH2of41sxy4Ci8aBYVoKZB4aIl9nAAh5phAB/TmU
9+XRaQP4P0ug0q7XoI7cz/VG2zvGJ4AFStT73Uk0DAsTOw5C1E/FPZ+4453k+XXG6Mc+9Edlyz1g
kLbWFQVeweoJy1Qzp8bNP+IGNMTCL4d7skJvQVtDKPG4p5whnWlSmAxddpd6vHFtfVECy0tmlv+S
EJrcLT+TUCBG/IeuSXVptff+isFxYvnnuhn4pIGuobrPDQUPOEEWqJwpN4vxYKGstZbJftv/oZqA
iGuptuHgJENrQO1WsB0BDUJHGq4UgoZDIVncWAJd7Qqn9T31exP/Ey+fkYN2k6Y7AwhySku120Eu
6cWt5Kw0wclGv1X2VJdQKGQfSBZkfHWNRtgSYl7NNmAeH/jhaNIK82Hj8SH68MKv1NcbQdbmiAjX
bSAeMcIczP6+kb6pXERE25oUFHJ7Sm1ZPsZ+ZUQv0zfdQFaA7UO9RVFbcKgktFOxRHT6chtSGiTn
sV+Cdw5pd/Prs7R5wPsh0gP8Ly5lX1vLSUzuI4wsrI/DsXX2C5QDx6ckFHxC/sNBxjsZfLBYWFI3
PKA8zV63kajeXm81USvUPZeskW7/4ZktpymFP22vlTNHtj5Qvh/XDpDlTzwKp2Xlcm9DMJpDN4nX
CvnlS86bvOWaVOkLaKVLMq0jXxEj5b+ZjbFQtESfsOYZ1hCPjWKIQtBsvcuuLC03Pgvq2PwGRtzy
L7hVVx/TFO3cdvnV2MK6VJHI9YEMW0Aw/7rNz8N6O4pp4JoljKWxJ+bQDuuLP9BesgdVfag1Ni55
kulRgNKo6h5YYNGsdR0fIBN+X+pLOcO6UDJSv+BXYvPtX/HPuVkBLLtitfXNULXUieo3f0NfGjgJ
tKLibaNRB9JjV0Jdy8SR1CPMN3QxKlZly8KHm4bj8RaRco5N6mS4QM3OF/3UiaE03xI9cvePLI1e
T1tj7bpPrE4gIDyJyaIMaCXhQ+716fPHJngTk/WZL2Zeeu/PLeaeMRj1f5i2SVu4A4lUJfX92nEQ
8WS28py3ABopiVbRbbPAxp+8lPwLDgi6i9UWgvip85mFnjwaeRxRfmeWzvhEmjE17nSENrqs6Lah
WTq2k+3PtPNab4vrR4KAR8IWZruX42GZGyLrq+HNdVfGj3WHIdQiEpJOATjLLz6Cze56pvfzkwKn
SIqkjMVJIH1WHuJUz0ODR+xtXfl98OJumqLe/LxN2uMxr9mC2aYAwFc7KGvskX/4nNXHPs8sByar
8tin4s3tuh8HtiIWU53NrMK21rwYzfJgj/9nMfsRGUyX9RNvKys43lmQh6o5u+zAGvXvbio7voT2
SIROkfkHE0kEZFXlz2Q5yOTW6OunImjpv6qPjafMpw3nFYeZphr5D6UfS/vHUcMhJFdIWMQ1hJ1Y
KXwzAO3OvVmsywloq8nNTv32Haok6WSrbVRqfS8kRElgXysgwjsUnqj0yY8Z8r8EDFCm9ojboG95
Sd3lapENEyphTXZ3/xLvjDUTo6XXLx1MTd7CY6ZA31I4rCU/+eJJEsqojFBuUKwZ9VJfy62PI+n6
EgpAChtTmGT0u78Cch/58MwKEFqfzd2OK3XsisFBDhxhHGe6D3gYpc8g+kCB/v63ZWffDDVbWKcM
6sjfwyhjct70IPfDskSHnl8/cI3ixiaPb6btNA7O9clRmmZoCbFsKCvpQH2wT4hXZfjhuG+6YGrw
BsNmcKWnsqi2DKLwCXGjiC6DytYVaa9Cgq+sFZd/kLoPvNbb+WA/upmPGrIDf8e2v/7gdNYUfU2X
jw1F/Kf1YxryOYQla4ruiWuEhZCUB2eqn+sipJ0f/1jMbBSo6TdQx1Fsy+DAdvvttDVFmecv9zDC
jo+jGD4RIU0HKjo6xST4tV21KAiTSKcPpTE86Tr2B2LFuLwPlU9PHvQFnWeOuvz4wt3ywZ+dRG9m
/0QCU1WhNlPj+yyFAEQ6wrx5uD1sU1MEx/s5SG0nNHWfShJSSMD8pDiHQkGzG5ujESJvyr+A5wHd
Bba16AInGxs2se91xIWSFmFvOJfSeYjCeUS4xsgzJsBuoFYua6PepYCV1chrN2sxqOtDnNEoG2Ky
M3QQ4skrcWlBTIb/DNEnLdceskpN2H/6mL9KSJWV/guJTwetgziF2/JR2Ei1GQB1x2ppFnZl5FOc
4nzTjohkqcRKgiSzLBFgCijCfTSoxHt+3FdEatX87jJp3UWC+iCFgAWhNNpnmt6K7GX8ZKmn4piE
opnly12IZFlItVYOPtGz8gBMfTAgc8Pazucp6vj6mhwNg4FPSsjo+C6G/x7bgqw6uBuJKN4F/Gx4
j2u2Zx11dQCC6X19Kmj7dquOWRapX+wuAV5OIbc1d4yEskBn+gciHgvIbr6e3L47nibDTf/NoR1O
WaP9nNqSOmbLfnVv5CmhygnnLp8nwos7HQptlolHj2IbIqJBKMWVAGeUPxf97e/OWNKeC4K/McYV
eWtakMTHTHwRf+MtK7SnTtt3ft1ZuiE1l5SNJEB4zGBX5eoXS/sO46W9dxdovTfCuKPp67xdIlZE
8jzFaV7i86KILsKhUb8IBYFJ9BxV4LzL7o7enAZ8kbliEM5wAG+pLHJ+BlkRlJ/Aku8LQ8q3wtnk
XhU+87uLVxDwCZ5mr9kaqxkQqGaz7UhnuwBoHE+PFn957EQydWS912rawN1i+ecMzIIGsxv6SgC0
+PSf4bhNhEgK8MOD34ApIV2TmKOjRaFYbJjfS+elzwwHlxVIu3Zhp7rsZ7Y9/8Ckz5UYOyquNsfm
PQRnhBuLC9w9bWmqMkoGfiDyFGYDxl/papZhP7PaoqGj7NgEGhAPqHMLthBFdHRFcB0VmTkEFGy7
UdkKTXRbkk0RiRHlQCAFixsZqadM52PBytcAgtpjziPwykHq7vsjz6bD+FP1y59wbhLr3hQU0Q5o
1Q+6WIBdKocy83E4aM3hQJgcasehgDTE/s8jdQk31+rhkU902gnqNhe2kaVFO3L/82CPpbRq2LSB
NeOfUdbv0EZWhi/ldSMZa8MCS3lo+nipPGOqttczvfSCjEGl+0R04ab37fP+48CCQly1TnsxqGRG
VQ912Vu7Peh84t3vj3jiLIRMXpk5WWGPv9T9HizHHfYtT+8d96XigA2msZPCwNYYW5WV+TGtX7QA
YZ7AMcCmAh6ZDtfiDz9DDj42PBzekgD8S2TZjaF1vDSMdQlMqI7bm2HRb81vutFvcG4cQjNw8mtV
TmeVbizzFX3ES794nNu7GXgtq3frAW7UhdTx1h+W8S+CjRkQmWayZNq8utN2qWwjl33e36KcbkXr
sy9wLgx2GIzXqS3wSG7Waw7nk7+oxrcoyVPVNk6NHWWU9hijH6rkWkUx+wzFFdS8NbgFq0bzDW0R
oVqYM8ShRkmMlz15AUcUVKXneibR4gbS1jXJmDZLZfaxPjLtuOGuvP1t+FbgROz7vIv1/cnJ4AoJ
bHTLuG21UX2mYCoVrqeZ6k7xTRgBVXeb8AEgIxjN0Jxp1My2ql0Kdi4is9qFqeutgmcY1esBK76b
+h4fp8hzZPv3OI2KapOgtjFAdbUDPBSL1oIp9ER7GmlVpk0zaiZbdx86vKZXRzswnVL7/44Eho/2
hVYCUzzKOK6IaDrlgScE3eZnJx2pkfIK/BIC705ZXgFY0Oeduk3/FkjkLCcPwiMzj1/eXWlR6880
+eUiI6xxWSRIHHysFVitvqG+wXZDQ0KzNgP3owsyi7DOTjAjhqiuG36vTK5pz/gKA2z23AnegCIM
ndAjcn2zTL3GCW9w3oP6VAzQeo/Rb2DDRf1TPcJcJGRKJpON7w64RIVUDqhQtCG4/WgE0ZBSDP/b
Fw4c/c4b8GsFfmBdu+AO0GcYx2QCpt5KV6ijBKGdjnGZM/eujufxWDkdXzerfQ/Jjl6k0fAyiJex
bCJyzw+oITsN7NVpWHmhaFh/qZ5j8dFiSz6vD/rUl2INWkvqriRpvA7ZgBmHDdyYBX51hKxf5OTJ
WKcy5ZUdXrbMguO+C5MIMBahdi9fCVsuXtMMX3x3GxE4d0dzn8i17gGu5UPOKZm6XG4YmFup3IYm
LynbeQa4Fwvo3dgkeD6XaADOVqFpso4l7dPQpnRKBHSDtojbgGmfmx1xUOevg3+s0gMsXzHKw6ur
JzRGJInTqYLkmg5XbrsmNTLHA2oEuQ8njSgbvpKcKYa0lQslZpIiT28bDaqJlOuNsjDJ1pqr5/k5
MjDrj4i1oHjvVAePL1UcBUZIM3IpoaJemtQEuP9L5St7v8LAuQlNgmO4JfuIPD6JGS1LZDZWTWXH
qmBHufkq+MqaZIIWgbt1D4xGKll1nQ2ifp9CdNvqr8G7nvmQhAMsg2FiVwu4AejITMAgJoEn7ekF
JpXUipTwc2jAKKval+838o/JzTZfjFarOUrfdfoO08TF576eIdk6ZHWfqfalPKZA/jzZgGFcdkK0
I8F7XkhvW90nET3lipAh4ABd3PgeAmMZhqsmmt78qBuTRRWytqeRULKwrrbQDj1irECmvDg+bieh
thzw9QAFnq6pCY5b6GA+bJxIXmt7vZHsb4iIw74Hmo1cMZWWllWbVaXIOcrZcMyajqHDbWDX2/wR
m9dGZTAC06siO1sJmzJ5MhtM55XsWMbWUNOO8RgTIhbK9gl8sGf4ZDL/uoHWLma6ZJoK5KTd4w/p
U2bwPYkDPCBFls4oxz1+1y30Pnj4kAJlBFe9HoVxmyM02iJlGrKudPdViHto6me0ai0PdbBPZext
vRhOiavxmG/sxBTVLaq0pnY4HiQTYT5gq3qdizEUQGQoe4KxtFdcKaRqDIe5y7hKenED/PmBJIg6
dxAfyfUnvmfscjMwlJrMEgpgQZGcnSyrz74oaYuGwbnQq27CPC+kbN8o5/yJRMSQLynpzWACbWgQ
WFlyOvsdf+GYbxSkSzZv5BmiQRwgfQwKKhVNYfv1zlh6PCW9oXoAu5FND3b+08icrJ7RIlWu48mX
JlovfGLpwkcsGIsTY31yQABh8xizkkpuM/ngoS6EH0kbkrgCtY5c3NbCxmt5D3tgFGMDBpYJp163
+ClVvDxP297/KpxCkbQlGKRi4+TsEuEO5h6v0ep01a91JQF7XQwufYKcbHaRr5C81MNanMYcRg2r
KOVDBTChQS71EqRTfrDq5H7EgGKxyxH5VsBGXoxaMc2Ejy6mta0slD2+G/N6ulGtQck2aiNyWfCh
Ja+IEJGFEdzdm+i2OT3/mdrRXnhhi/MN1TvSxi0B7de6uZEk84KkmpI08fq7NdCH61+N91QkZnLu
M1urkTZiJzCqTlsT0XgPavpv+lICR5dBPibr3Z/eLGguGlR1XFyO/5Mba1AsUablJV6tHT+TaHb5
t9sQd7uVmBLKcew3k1lgPNzfCBqH8LA9BrSgiPMmPAWy7liK4esS1iuqyL/oca4fbvSbHMTDOAhP
YLxxgFRFWypfaSEfLop9vlarW5CY3A7h3PTwewnVIrh68vh6I96fX99O0YG3Wb/jCodg6ve5OmAq
L9PyOVFhNLnfFNLRr4L5FBgUjY50VtTdjYA1cYdtsbpyLwAVW9elbfy0XCufiH6uYUYdUzYhkQHe
l80MzDua1fjfhKi6PrukKXXgb+eqSMB+sYWH12KYQdLToEm7vJLPvhRtZBmGKp46/3qTO+xLGXVI
T6Nd5MfwA6xEvR4OMhlweBusqFE6w5YRGYmy1v0AkDYgmnBkXiMRw9po1w0rT1YG0zBlEURzL4W3
NbIRdB+CLA1NmkxJqk09YOzJhqn6GM05taHkZkkJSHAKPvc9Bw/QGoU/Hx0FGHEsvS8NMyocNo3r
xF4H5q3UETF7gQ/Er+G73r6pflmcyB/QLq7HisM/QO9m5M8TKLLMLmzkexQNqBS2IANWaWiucSVP
VTXTu+YRYP/wkNtlz5cSq0F58++dAFUeDFULuXg0j669igBlXiltTrzG2VR4f+aEqh2lZJAhvHNS
BWRSWZsrv7ggoJRzwDynebSwZlgu6OfG2HeKBtC1ONbaJaSSf4vMwhd37W0WiQJlFfLGPKhhlFU7
apNKS0q7WRKLdyLlMORxPmkmzMRcdCuWHQ19sNf2eG0op1G28T6UKTVGINghmSHhBOryGW9davHA
meb+mtKw0IVmG3hhBACqBElK7zm1yI181HnOUdMabkCpYGVOIGKuFO3WPRVpxHgHWNjgP8igIfNV
qXJ4zziF/ZgSWv8s4ELCfcwF6toqm6ikbb5ecfIT1ibsvI617UAVzU3/pqGClNjw+wLnCjVfx4/M
UEMuKnZp+KKuLR/FfmSZ2GJ8/Lj2GieFpWcWjjPkckBOh72y1qtdEi+woIiSUKLdS3VJ06UV6l+U
UjpcPKI5QX2cS5PB3PV0RYvMaRgzKBWoJ1QE8xARpKYdDX8K4oNX0TYio169vdnT87zdsJd4WtrN
GwjAuwCJ7ttpYfy2UgZsb3wZpkNMcElyK7ZrW9QYZNFVg+zAhEJmoZ2ucIV1TwiZbBkDNsUYMsvA
xIM5FhxjN61MAOGp0qGGa3pvsutyJn2LzvM3GDFpQUxjZciWX2LQ2NdzCDN4zKmyBU5zYAof0I+m
FkzKqvtVweAme28CzUHgXv+T8fiKBvLjCnvyEs5CYx/q/JxaNNmShDQnqZOKaGqRUFRKqU+VGxLw
sWnKAQFykLk+oinfo2Go7E+6AcHToblaGzw6DbGXnCr4GloEfOPhqHG7b2z2BFvgEtHb1PHHL585
vrgQos+YGd6ThMSjLbeHuf6YMx5/R9SCdGzoxmeOLm4/lRJgfnuRqz5ddE6U4Qqet8cEzmW+ZYmg
RXSw9ZQDZwzHszvOXUKdY9fSErJ6eXEISJnrxLujKB9OeivY5w1yPuJNu36wvC0QI3oXxUlRvFrM
pj3UkrfOYH97EBaQmAN09BArLv0bmuZrJ/JnrMFTT7/+RpSF0cEaKnEDE7GHAL2URwCwIrputo1i
qNbFpWLIYbMXwIZRKDbhNG5jk01o0D5boIOLCfIIis6nZiPBX8pdcUEJutxzEsb7qxUcdmpf9Fxq
f+eTsUqDgqpQkz8sC7us7LeJ6Jw0dJitvRa0htEbSfVlUoqTaW/Hh5YUHVkKUYVW030LTO5AX+uv
YkjIFa5n3Db2gLTRc7Ce40JxJDIQqghdqKhIr8jYkEG+r3SOifhBpWE5aoEA8qJZuz+41RnntS/l
wKk+JBDeTc59h5THajbqcQAfzbcvo3i4KHUNE6R/oOOroN9rdQA41xLrzsdvUGr9FFB3UdWSIwRE
Kvh1GNURBhr/AH+iAsWKNJVztOP1blcqdSVCTwvLbz96bnhEhGq2n9n15RI8godkT0lvMn6rOpbV
RslF9X7xoe/XmUA2kU2kko3U8/NDSndlppScVpqgDqHxdHZueQXZs51P3fstfgvZVmkMZ6DDdV9P
Y3aXweVtQXDTfNlcvFkCdVjIBpDEfBHeHkWZiKR5yRefryK3PJxnBHkpud+Vh421OYK7HHCyr0M7
wcSLBpWVMjsIQIaOKrugO5fKM8tKMIyIb6RGoF/Qx2AsJPBRv2sX0k5rHKMWFPFkdtS6UhavZWc6
CODyQggMNq9k2cfyl6BAQxsFd83m2qaCETDbzcz14Wk20X7GhTlfMuQCaZaJAfZgE5dloSGJQzYZ
pVtMkYN386BgG2H8XmiWH3Z7Y5OIiH9vgc7iMpso0f1zyfN/vVuPplMEgT+EqTe1v55dA+F55QuI
VfKo6OagSGOi2efHjZr1fKdzJtMsfqUYM8BYudWSRtePwdfUH9+f1WyWmmcwWql86X0beiXkxmpS
38H+hXwNjMRLCg6cguuzOOhVfqod1hMiAJdD+5kH9ycXKB6iUewY7qbD+tJy2mVdxGXnUZlWzrj2
/ccJXayUAD+efiJ7dKx3DqwqG6a+bfHZ+7VnOk4VBNKqnFXJ+E0P3nLxmNg5oX8dhk73qBmlvyvN
2ORckp4KRPb77wOAyu04S1NMpXgFicFlIVQNGcLhzpYX/vA/ucS5j34e4YgkZW1aOmb+1fqc60xy
E27M4HfGGOn6WBTth7G56L8HYcJAJWHFEf5l/Iar/JSSc6JXlzpd0L6f5Go1Xqr2rnfx9RFeicgK
IaJ/VE2Gv7pRXXWWNB+KdhSQLKBvrrQj+TgRAdvINOWjRzoT537+7pSJLbSK98SsYoU+X2iOZHSK
FMI1HrCwGrm/pyzQFrJrKj18m+C8TDrpGwwfTwSJDsJHkYHE4DqwuiJF3YLDJngUKwMkrXREKDBR
GP3dCzOYmWIEHysMGMiQZJtkxTNb1+D0xJesmv/5Z+T6/kB5/GA4FMJxsIZLgai4D70BphpbiCnd
wfPFP8n7aK9SNC7FQQp8Btg7amgnnxm7/LfWYUj9kmylJ3xo6AGFk0NyDVcQu7B/letZLaDdZbyl
zDHj1NB3Yexluav+aH3of6Y684SH+88Z2J5DVezRK5PmOcMvULKJxpfe4u834Gfzk4R0GBYX2ACK
Idd2CpeiX3hR9ZGQ0KJQ3fdqXcHGOoV6OeWfmgD5JyYJyvlbGeKV764Xbql/1ZCRJCI2fLv+Jtzz
8eQqemikWKjCLqJq3NavzCn4B+rrd0ciX6I4v+tp4SxVdGtanPpVYDx9r5SCczsKec9SRH8GP7q+
r2E6kVThgVTZhOwj2P+i+EGEgLQiDDhYkRi24YqtCuNXMhn+znYjYbjFeecvhoucLiKj0EiOTfT+
+E2lwSKvcvXCHsgw6zgfHQOojISrEsKale+nyZlndH9KVOFEY+IFvHMpnVwJtgs0ZM2021SlQzf2
Guqff3TY1GB34ag=
`protect end_protected
