`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xhdmvpu4Jx9ulRYK1bms067P6bkyvNmKsv4RYuGPBcntIT8Tv1OXHx9d+oma+1332EirWw6dfB4g
xXKY+8ulCQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BAfl/GudGL9Li3O15MBaKBn9bId2TiruFEmoazneGbf/D6BfZ8a83S4BWNm+JlYIBB0LqvqYftHL
v+J843jA6P0FrMu8Q9rPf2t3RaO5TKce0JYrffzz6G+RgYOFVCS08zNPYYoMexzkRcN9XarsTSZL
y93eGAW4tX1W1y7DvCo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Xx6r/Bb3xF+5/QAYxc1h4dAQRVevozVWN5Yo77uoyrqmxwHl8cBBiMbCAj+GS+H36JgHMjxbuG3h
dYlOfB/ZwHBdfsfxfgCCrC08XdPrFiYkHH/cMFgAaEi3jod9YtnusuaqlSckyHGBEH2qp23YY4OG
UF2+T8KlU+7D1UmPSjr5rOuo3ffX0ia9EkeZRF/F9s3njfsto81l/QAO/A30crUK35lSY2oRgFra
Cpp06FlHEApIyLZ++xmxttWfuTdjH0Dgc1sE2F8jtP7nCf84irk/ZMN8yeeF5zKo6nvdpgwQbJL7
SAgvcHjHGxieHnuVrsBZvHesSmLxGRaj9xAXlg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Se+g37Xd/w2oyxNF3kBbjhMAIoorO27ObzGbOxBCQmD2SkPtk728J7zsET5IK5jc31p4NEh4LEZV
vbHFcP60MSQlQf8HA3Vi4+oaiQ9yghe3cYunmdx1xC/BGDyTNgFqDrtKrwGyHiwYLr/Eo/QKTB7e
+LfSZYtydBT4irW1vCc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h+UC8NP62XnpQpV3p1hp4ojOn6spTMjTLGw2+8Up//qJlg2R2EoYWeFS/02NDAyoVMQmK1bXojzS
yMpp0tjPoHshKeSjIHQcs8KMhsvuRbd/NrJ89NIW4dRpNqvXpjpZincbLtsIbmFBpE5TKCgCfone
JJYB1Ns63hevEXSs5JqDbkLQOZ+qRb5csolUj7+yHU1Fj/VETN6jzQhSHUW64Ewq2uaqg6XjMgQ/
27jRoWJrJG/wmEKoK73VwWW0BEk9H59DSwMcEEbZ0s31fuBOpYDtWbwFTQ3vU6Lz00t0TbPSFlTs
0fttTMI8WOrdcuVsXb2+ULwYklkOkM75AfOOAQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40032)
`protect data_block
eEe4YsskQmU6HvOroUgzSYvKEBd9H6S0bP4aWbYWINkH54QV1A6z6VqlQsxlpzNhzDgR6uSMZNpS
xfGs+vpmvikrH8eiHjKfxUZ4NyuYudYSncVETpJD5URhCP91P1pBxYvSGyjXn4jqIA0orxYBQbFK
m5hlpKaIFGzFGgr16WlRMTOdp/+ySwHg6qjfVtLxBnw2lfCvjpLPtmx7unFRruaguAHQKKoWbqMe
K6PgiZXodbCSz2cNZutivJMYsJ0aWfwxb++vkDc4wG8xKeEZxIL7cDPD/VVBz1kEu4Vil0aJfOjm
FUsVGob7CB0iCE1zRxf1qT5xu+uBXexVboOFdUdbmBT/40vptvFGcOLw2X2dT8hcsya2YJ/WfN3v
P3TDpOkxEGZhAGKtRpPCLmE+M83KfiA4G0VBNtHj/mkWIGPGRGBOcTlMDrXXRySadyIAbENTD2T8
XfamcEnZHPIfzPXjfH/osobU/JgX1aCQjcKLVkHwPQRxvLfA/XCdE21+Md2gShBB4RuAX1eGSij3
63lPNKkQ4hFugGGBSilmo1mfV/NDJuL8sxnO7UBhZgYI/ttXewafK27PFKTnoFzECdkp3r0PJKLW
zwNIsVtqrEtWjg4I8Cmz3888BFuk9bvQ0AW1fem5oQWIo/G0JRMBh3hisqjqsS9yvGv/n4gZX1c/
FBw+T6AwoXztNDsYuJUXvjOBT96XguEx8QePpWPQwilIo3qV/oy0byKX55cnP9nh40qxH4NDAjR3
OQO9ujX025kl3TetRcEhyQnKr6Fc78cUMSnlU/UrgS3yQzNu1WNcOTaboZ4QC+MGzt0rw4AN7m68
30O+re/lwxeJnEYUARHTGOO30QoDrOV2AdsmABeEE9PJpQz9bf0wW/M9upXyOUTe4TdSPUxxS/Q9
5+/eXwGtltvdvHkAtEIcuHUR0/hCrjdKNgGNeYL+s+/03/sVsIXN0bznVMyAPbfg7g/w7HMdE7EV
SMxt4+zwnHCqCn9Ln5u5VHqfIURpxfLWaXb8ekgoSAtBUzCwQTMHzhZ0yqVOE/Qcgf9j9tiUZio5
d5Qrh3+nQKxvdkl7NQ2HkMKz1cKxBnNKRW9K+h/bJxToHcC6C4RS5JEHUNAkFWXNiWo+UYcnrx4t
kNZKPfG+WVn59Y/QubbORXhm2/QgL1gAvxI+pPH5ZvUKTDnylXvQK6DMujnFHUGvvXT8NLZFQ6y2
GqqoRNbHzsXU7dHSFNCJ+yts8V6YegBxlfiamUOQX7uh5GcsZa/E+BNlI0+GIo4bRmoCo1p2uym7
MQdSAhDrDDvVHYXI6McRtHM1gg6lQwd1xaMlxjv4lQy/C3GExzsDxARcAVcnoR/huLfmo36XptEW
wILURwNPtIl6EX6ZjmuyHvESnbHOiLo9VcTEch72g5OgTGxihYu8r1UqhSOWU8vqEx29IRju14X4
yB0gi0cnxV9b2dSwH48cF6MDCFUtvFaPFmY2x0WmwUrL5xRjASty5IZOVEnTFBk0fhm7wlJhk4ar
eIBKYjW3ZgEGKz8CNMoEWf6pNihCatCKxRQf3ym9czLsjxW1moxjj91yWJzA5IgJ3erG05EWpffq
1egCmipq4G/U+F1+Q2xcZ9RAZO0I/iZ76ITt6mGfVCEy5pvhEIqIbwe1fiqsRpzX3Yg07n3wzc7n
Gvh1Z9XfgmVfoxmeojQ2eLVcxrllNRZFX2QW7w6RqhNpZY1IQg4wFbEEBiRdrOV6mLlLZ5Pl255W
ZIcFNCqGL1t6z/TxJq/+bpWMz+BL5yZUFJO7M79V+rXG3FmjRIeKvdzhwONgJCeHPCfbhkXyb58j
DhlihlSMaMVowsY1F2+qz1l7Kh30+AvTmPfBtLmot4RKa54JV23U6+50sGEADcft90mgerAk+RfQ
xiM5FRsic1F/YyKmsmb4Xlh5N0MKnGTgkmHfzWCpmDyO7J6RWmDosOcqV/h8bF8Oxx3wExqCOzFK
1UXVN0ACCNHga3PFMnzILOZAZEnmxkhST5wNKz2IhJJqSOkokwXFZySyjtBllXI8diRvY0hgTGN0
epicMZAFTZcjP7Xk/K1ZD1yjYSZddlspQQ2WvNIZ9+JsVsx9Rs4TBVCfcAMmclp2rFH6MhIuqPjN
8YrWVUMNDP1Xyrgf7mBqeNXfvWaZotyG1LnbF2yh5e9lyI9kyF+VCGJkUM3XiGd5DEXmtVkbFXEe
C8UpYTuVFl/XJeteyIETCDZqRk2N9Vq+A7B8ZeDImzKXB6eQnaqQ7GyZA3Mf22s/wfy1rcUq3XA4
MtVFVy88wO9kHH7MBdPDp9KUiflXZar6lr0WxXBmhgXRNJSe/f6S9ohlelm+kdbATF8KSK1xAj1v
xEOYjWfXgb5TQY9MPoexeHAWS08onDir8orGHuhiNTzRmcJzP6c/506phn0JQXAqReNFF0x2mEDD
+eboE7sBSzBCDQU+eaAmmpxHcYJ+D2B+Iq0Felm73rqoHvi9tR2bVayh2RpK/T2m55J3kTVl6K3x
2v+Hch74DjXnL31R45tc9eYf/tsh0K2CjoBYeiJDjjzL1YctOIkuYBZoOTdRb1+/IxF+R5ljqPuA
sCjr8B82I1D0rZpc/mGYHVexmTXG7+/se7qZ2RX0LMq3/8J6iLeR6zmLZRn1k9FU9Ky0xgW/Onje
VM3ujhS6iWT+od+lu8X5WWu4nDjqM+4O3MS7XiPV6DsLxGC5SW2YiOEIPlV2rFvOCryqnP5H8Hec
jkEwjq+s2fYqdmpQQ0V4KFd2qykUa4PmuOetN4o1vNQvl7kziyM8WzZgOaUlLgk8ZkWdJY3hMcyq
urZqtVzNAiNh6eUqcIaGTQZmw6QXoDKqa7kKT3aCWayXTVdngbTsUcAoHBn0Aru7XW844JSA3GU7
U7lnUELVMToyVOdUMRqwRDuxWgzJon+Vx5JhGKX8fgmbSvPFmzZzgmTZN04+GCouT+pXxwNvtPsH
6gsUWNArUpzHb9mp00rByuaiHOaXOxA2Lk74kn5/Vg1PoHK4Ld69GpkdybEYjnRBD8HrUA5WvkBQ
dKjCMC0D27YJdJCa3qSYm3XgLzd9MOgsDhjNcXsOre6i89alkHiVjGT390QYQQxBWlOoshGJKd3H
nNXBcx+72Xd9H4tO6wLTFCy+JEAM89R4V57d4G2vQxgYsQDLZAhKisSTumvNy/41J/iCXSQYCWiU
b2GUUw1g+7SgzzPjsvCFDl+72scYiL/fbzPOgn5wLhAULFOrKB+ft4fV2cIEd9+JrBXfbK3Ba3eo
h6unKFO9k30GFXg1H0r2fPbx2Kd9k9QyeUv/WNOrDC18ITedRC/0lxOmUrNZCpcIu0/K/fVcpiv8
6NTGTpf3QXhHFa263hjgLd63dRsyUxDBvqjnFOiPTEtRA0KlMhh8GiFJxbDIvDXYBglKLHB+Abf9
1uiKPJm/7qa/O1zScCJAo/al7wLnFgvpRt8UkdXKlV2OkWpZbG231FBCOLSq2kiKvc4YLxrWPU77
31vj6L9ju1N6MZTGYl8uhvAW7og5h4JsVtckgKhc3IgSyJ/4iBFauIU8k0gCpsOzOew+hkOGwAX6
xWdduf2Vtqu4D5+OUCsi6STOFQVd/DqDDOmLGvg8ACoy6igoK418nSxxN9lD5bP5ifCYgcDIdHVk
Rdlx5ZxOzb4Tj62UCW7+uic4GGBRCLjeehv05xsWqRygvg6mTUMVTdGaOliWTQ+b3aQe6gJuUKyd
Z8S2yBXeWyITJxmKqsqArZGr3qYJhSoV3nEqfsXSnieKbbs8uj6KwR8XV0TIPgBSuYshyILg3ho7
dhZEkEsGjpz6DD3KxteZ8fMwUGexhXLDGWfet+iXgnZRFBmBJ6zEU4C7yeQ3/aq3Su/8aa5cQrif
2zkOzM6ITZmzfnPdeG1y20wxzko3vyvILtsBWl07W4gWVJhZtdJ7kRAqEcbxWNgH1URjoHeF7JxP
sDuhS9mcttcNRWWglE+/hONtebSRNG4FN+ULXcbfGAQeD1ypDwpsYHBeXph3AYYhR9nwKM2gkTUP
5fYOL4oc/RdwP8HhWjspfCyCDx1bKhRANOhftu0qTvSKwCEA3fGJBEU0s+6xYdEuUlyjlKLOLTQi
aYuB3gZw+u0+kn9LSMS52CSwRKDBhNyoGP+eGns38XSn9bXs/7sWUREPO6U8Syo2EUjTZOSySeHm
2IJE9QW4b7YDzgr3qnqu/hSzSpVWMRdAGhgCANh0zJhFY3oNrs4Je6zxJ86ObzRdkX1U37Q4tCXB
pLElo8CL8CoEYgALZ2tc5Rn0/hEzL34MDIbVoGgOAc5T4vfauW4lVSnyHRubxD7rParMYZ8kZA0G
ImsPwJtDyrmSkX0N7Uz2ebV9O8lALOuewIunS89HDyK4QVAlWTZrVMaGH3YrEKpXlaIv8mRwO2jY
zbvQJ5Y4IO+VbK2PzTwtsKex0ObEhSEMqSGuX/vOc986Zcqh+XUD+MDQ4vTe4xXOLgyDriUC6kWg
vClsKthUuyo2wq9FpXxLqACWXEHmgdwgOkMj0GnPSJ6bgMtQHi4DdD7WC0DsK/cCouC3lA21Lf0v
srMng7PRF0bEXC9aX5UGeZifLan82AIz+pyYhnASkEoCmQBJNw26gsCfWC5OyDTUnLp9k9puau++
7WEBGHk26QjvBbyfdKXimQeNKhGxu2xDurT8WZ9pWQ1ko5ToHZrhurzeR6gPyJn24AL/EqKZmfCi
l0rlZKqVfpi+s0MbEZvZq0Nf1ZIQv/HsQmt205YPPgXGg2UHvBuMLqOzYxklor1PLpMaB/try2fI
cYqeBjc/DnIVDGNmINR52WhZx+rfoIMB85jNkm2ih7mRwTvLP0mpMRRB82Wj33+p7ghzLkcrBvxN
delocE8uISJutBhtloT7sl3SVVnMoUg12PLXLDEr7/vFtMOeLiWJHvxNuYdfXa5YhXny6/gtn1fn
DiuQ1va8X+h+D4RBABpPu4WKsFU0+i4iWJpfkahg7QqoDfGhWAaYXr1xHA5XVGB4nIViUS84X13B
zdK3dJCWkMpYRgX8rkwtm5vtew7/uMwlsVHicF1nahM/2ehWHJsn8BqSAkl03Ji2KL3TPYPe/odb
q4+GCibcZIWy96uLxM8ByX51O8Oz6fOABJPe3YUBEFJNQK7am/Bom2Ft4zpDf8sRDdowYJzrL8qX
6Y2THFmY7iMyLK3a8OfSblpM/68tBBNau/CtJUmJq0L+RCPmvocCZRcVJq8geXWFfZmoIc4m8Ta1
y9D+u6aNBgQh8nMioTM/JmGkcBWUhX7CMIIwycLJ9g2DZbQt7LSTg3uo+0onDaPJdDtH200jNvmP
wMeGKrecA7SemQ1ymcOKkyZxEtj238hYH+YZGnJgrnhX1Zop0UcYyUXxN5nADZVe6NyNyUPK+NRm
P0+9uEp6MxZEw68GJJ+ynMALwQ8lO96FBEDtUrBW8sXjJuLiCaeogtw6qNW1hX6y8IvD4hU6NYOR
rb+coEqry58+skqwCkbZ5CEqHrXLfSAA3Y0izQC0ZhgR5QaKwJ6T0Q18XXq5f8TEKa3ZMHlUER0U
YK0U9x3PMi7r6FFzL5U5LQa9zSiTZcTyJnrgYBZIdh3gvAm7pDmFiFaf+L+XrkHAMN/3oDTjmxB/
Fc7BYd5P2qFf3WwahO38ji8Oo9Nzp3mS37pMjJUXASWd3MVfnpq8VOmzIxTrOUzO+jXnFJmr+Upp
wHmtn+CqXBLp4XJsB0rrZv/6PvyCZfC61uu1A2c6AueHJ8sSwzkZzk1WkeI4VU7Pdx9Eu345MvLk
qrB3mnBirxFksQ+g9ts1AP9iLKq2LwSBaB4wxEAZtK0YHSgd70v3TWuD7yxQL8joAfxNbWYM8R1G
d26Gl3RBtIca9mESpI+7SJR22cNCN4f/CxS9zCobSkDBnCwmk1rA9Nnb+YvJ3ZWuMO1hZorrC3li
UGuvlx5SvHHf8epkItYVrMHsZxclhC7uCSB3d8zW5FDuNJKD0WcbjoNN7IOzyoAniQdOuuX69XYl
ID4wNYxszDsR9ufggCmC9w4GKjC2T1DQC46AghQ4jH7/PkIs4v1wQw5MYiBMm7PvqlibRAP4jPLt
FPzn+2meFX3hp2tZj8FixTgvL8lgO29v9DXardEmxl727ey9UppAcPTfi1ab1bIyBvUIdYjnC51n
0nnDlFHkqNYRJBI/dHiK67UrXbJvq4Xe/NBoGDe+8TmI74GMSPMygglv6Qsvf6+N9vEKeFBnrqbG
Mg1PUN0FzmtTsDRWu1ZSPAUdAg1dELQLbYsZTW/iDgFy9XsSzjU8TJVZtIsufznzIIFmEVLJH6Nw
FePt6ltBo4iabuwVs7Yw+kN5OoV14Fa3zfPFevB5ja5KA4sX/heGnvG/TpQI10xERfOV19k/P1mK
rbeKoNwn+OTiBA14yb5wu9tDTBgZTs1rroEvLxyGCoI28P2Ljae9iHGzcMCt1Z3oIsNszvEi/z0i
s9uId1sXbES5BeNSQ05s6zXopkAlFQY2xCTbV+kn5A5P0MU+8Wpe2OamP7kfZstFCMAWeqSe5cWn
L9NarxxJ+11zT9fUIyKg9xXamaH9uFAATbSxWGCleDY6xknSxQc+J6p8obGIHE2JI+PYUzRRScX7
nRJtRzIEuTiAWQIU5SA8Cvpvt8lPdirGnMjX7+UwaXbcnPiUPaWFe7ERxWUAzrCmj2SWR9IHECwK
T1mI5HKAzGcPcPfkA9XgnspC4PM346XOdme7dv3prHkW7BizMF5+yyzTQ97z28sJUimgpa4ejG1R
Qv+zCTKonW7gvAIOkV6G8t7lQXWezR6TFv4G4pwjxsXAWl3r2lJWe0cFpZK3ex1va3wkFIOn/HAa
R8zhCM/R1sYUmTkGrTrSQeFZwuWtkra5RNbs3Bkl86vg/aJ/tYG2BatVsB2qMsL8Q8LTesL/vjJc
It60QuaR628SpwvNdAjrzDy1K9iQ/KHPWUKrZ+lKKwBWWwayIxVFw/F6YsKunLiJapMXFZAzdmjb
NumGOzIk3DeChiL46jSrxILOefD26EabQGjyakIEE4wfKG5PMZONDX8SMubbVjkG8MLNrOGXQ9qV
PpQodkcdDRngdquTH8/8ihbTAS+jfR4zVNeGo0xADvk1yAmYs2lpXk5VqlgkoiGvTCSx+j3Nivkr
Jwrpm6r77yRVTcWxhhvDEmoM8AExVpHv4x82x63J/94A/cA4XBY3jaRYo0kGmTflpy8QLSCtMLcN
msHvJRPNs2z+nDh/IYJ+mT5fsGzvhtBAvesEeEvUR1I1nl4a7VUYa+LE4lSUJZzyTQ+j1tWSDULK
ajY3GU7Jnk3njHO3svZbqazSFCP6ubfbD7XRMaqxppne4NDKo6HgScc069r0spf2mfDr7yDuydNo
LXMf6H2oU9n6QCStQHNSQLQeq2XvuUoUMqcpt11rSwBhQMwGiNk3xfKVowWTK9Pj/Uq9Pra9AjW1
PMVBIxUNa95OHWKU2m53ILFzxrAH1PrUw1Si/y4TvvWrMhjhiOlS+Rz1XNp3h+dd0maesyMgmp21
0PhYuR7bvseHNArljVoSJFugNkosWm0SSShQ4Z7Bk+MrUFPCjMLce6DgSHojtGy1Bsw4CRrX9E4X
n8f3bHTQUx9TNSsPayyP4hmUzYuzcyBKJPM6mPM9UWcI6IRX+C2sjoyVqAcp/LtVd9rT+Prv6URd
8mTBb0FdcaWQxJhwJJEe7GubVjjeSrH7LVzNzc7ZKZiOg8fX/ctwS5Pd9c2V1d1Hp5/Kxd/juh8j
IFloSdCag5g+uUTlWiiTWy0ER52xUgL5C6dQYJXYov8FM+gw1esnWRTGyyR68WXwTJPpSME55gQr
f0bAk0K6F3s5dPHI8qGDMzMYBpS6h5ggiPKyz6XCzeuP6n0ei9tB6jYo0fGbD74b+Mf7rawJFoV+
5FgRf+BphsTTzAXUM9LW5a2b5SYMOMuTQtlTp96P0CqtYYWfKJNSV4OcyVe9J7OCpfGCoKE41WMT
/dZT/Oo3ECy5VDy6PkVmVXwYxA5mmbSw1dZ4aDkB8xCn1MEDHqccOVN76PNpcuUCTaxCWk380f5g
kWPwjYxcIjDz+96L47w95nz91FOi3nozZwAMZGtTBaYrXRZ6zyozchDjiE4cITs1mx4rzOt/eli6
Dk3kc8yfg7oS6cMLU6qcDzwm2reviUnRfjtIuvjVuEfiWJoqsNSy/LJJ1+j3CTpT1aG43c4OQkv7
sfhcPoejM/sdYcvPH5aZOxvVs01g+Wt1dhJ0G2VlDRBrpRUOYfs5heQJ+qwDn+9fgdyAg3DKuafG
gkNHeOQNSQ5D0o1vHF7iopSzuFmDVEv9LlSTg5DFgJf6yd2b8gL9TP1IqnQSrIr+uIukNO6KoaFN
ekkRckwuBmSvKQZdeauPzRliZ6d2FxB//TP7CzbS1OkNMK+xgT30+anH9NwAmExZuNyqcq7ddRYR
K+ptZsn8/RbE0I+Dv++zGvik0iMwQaFL/eOHHXx+WMhe361IBdXC6eiURo3DVU7uxSq4C+bkKTSo
S4wBX6HWC6rECm8T8i/Vo78SUOzPi1aBcjge3O4ahELLBBKaPdsywh2pKAYb57EBhSQQl2nN+Fdb
Yj45AmHkZI3M6n6B46IrGR05GI+KQtS9hhTpzN4m2tfTF04U3bWhDZ0BIc3BBCzKh+gRsEkInuQ/
yyFxgu+zdHpM3HyGdSVfU1ZivEmVCnw8Al4qboAoWPJSVefKPAzJnDbcfnMKW8tPG1rgUUVQTPH8
t1uBVNsOLjKibeh0IcqqewkxMHoGuDoKhzQdEYMtZrlEaENFvuEN920EUkOPuny/SM41M1qils4S
V54MPHUq40uxQ4BcfSATvEBaFhEO4iGk4IPzi6pzNqHGviRXBWdKIRpBWiVLDXUfaHos7mPuUDuY
QDZ6DvoR23NJf/E8329BuHOEJtuJTdghZs2CKJJgOdrUjW9kqyQI70ncnDYaC0fRqKJ6CpvS4kyn
BnXOzhbosPi2RJXjM7aChGWRUQNBpYOUKLq6qSqRXsCkqZmwEFspfhfZuFZRc3ChpQvI9XyOoyRW
Mngc05YuhUUA+V+xImb9gMKkwuxGedMzS46OXtbiTjsloYghilbn3fcdENsTEPtxBaJuYlKE78QK
mKPCOZxMHNsVvMUnEG09NAY861KGo+oep8UZlG7OPo0cZZPP9Jn+OauvtfRI9XFXGuMvIVrL89/5
Jtk0Ncu2hqaiZgUDD6b6bXnVxKPvGCRFEhOYjuiUoAZiogJaYbQ/nleERejL73BaCS/m/vDjKP4l
osZfTIQ4CNA53noDJZKxm77rJxRISRVZ6JOQN4nePSbz1bYRDZJJ3Ik9aFlummMnYDmbnVHzVPCW
RyyNsZKLOlJXCJGy7cHyAYlPpGlf6tHE2eVCKo4cftZ3342BhiCbx/f8eWELdL3wVr4FIbjRYWu5
kQxWa3QnIKqDVzPHKuMtc5LXacY4TxwkvzP9moVFoz8qrc40GlTWgBWjhmQVHUmqjUa/AjNKsJIs
HFRHdRaZBLPX/qrN0GxPyXTw/qvHaWkjlAMm56fIfW7/6T5Zx/Te97qOU9qzulNH4uJorslt/saZ
oFkDatx5jONhcoSgpAXHZlyxEvyv8nwFeqyMVOawAGMqpe1ec83v4eM54xFr/F6vREvjMRmYxzST
PA1iOo+ZYP4h6gCoeNpqLVjQyARTEFyY/nr5EahBbd1wKukEhDNTHgTfbeFNsg1VbivMieBmLy5V
n1iKUH80Sj4sWkaUsQWyY2FtUKjGK2eWwgmLR0NO8nlIn9jrdV8ki85l0d+GBBI928CZhVwhlKYX
coAMuCQedrd6snnY3zHmMbObdckHLpW7u/UEnEw1SHBU8edOWYtbswRf+7qOeWZUVL6UJAnbSg0k
TucpiRPE5dfJdGWY474LeiEqLxFIQwzj7m8tQAwE/8ZeyLBGtIUPkCZroA+jfidfGo/gzUzRJjSh
FLS9ixrv4rXfiS5U+4qfBptGCMAIUFv1FIxkMaOdlr27po4apSINmTFRzx6/DTACgtdpJNSJ4MuY
nTjAOdZTmTg8FA1cO0Or/DzDS5S24hButv+qV+loenzy0CWxNS4aauzvI2BJ7Er4pi3w9YL657zX
nteCEdSUSKnP5ulA4yKDrONrbS70is783xOQZF7J/0pogjFAwecM9VjPjcNKZWs1ad44iVz59Y5c
vmlNcUcv5R/dNniufx26UB3CIqcyZasSqCpFOoZOI6Fa295vmN499BoWHz+TRt4zEA3skU7SDrC9
n0b5lNyJwndFdD5OSP24OIYnvoKo+1Cl/ZBVIETxxf8YDatJEePFeytShY9uWhMVeXhxB/vvXv89
BuUuN9mEBPtNqHbO2tqjQJYQc8bHE59ni+IAaIFHOChTLnzKYjQ3RPpQR6/0dNtZzcg0ERCblpuC
xkmJq+GjfTNtjhFkPp/b651uWkfJVLSaOluWfZH59X2igiMeOy4xB9nN4Ss0lvqJO6M4gnwJKcJp
VnN56mR7taxxwPlb2oUMs3pOKOU6/mVrd8TzvfTkCDtg1vDjMkKYj067IDn6onqKgZkILoCfYekC
SVe8KWYrGOB7Jxb7qKgQ1VH6OtAhoGkumyFX0j1svqrIsFHeFOKxcYzDYNuyd7Lu4Grcrm741FC5
PCnJD/q4pDvGrCzBoLfUeVIYYK+EHSWolCxHU2K6P5r9Zuvzx69YA8tjfF1Dm6kLqrEhhhKYj8eW
nVDEgQFCwP+I25sQsIxTgluzAV+e904h/uYPFXIbq0qkBsOOJCsXCF0DOLePpVxmkXt3Ag2yqASd
H07+7uC4sOFRzomXFF0S/gI7YhLz8U092LiBm3LfICQuXchG8Pu25z2QcqxETjTTtU/Rj0jWmzwO
EkqqRmY5mC6WiYCVYpfYm9Ou93+AxkVgDDr4BRB04ARaGed6ZIgffKD13QqCtznQhxRcM04HjncV
S0TVSY2I4daEBU2rQGqr5dXNcKWxQuBK6PvVjHUEwVZa2q7FdDVgGO+xJApfDSo3R58mrPkuxkxp
3AjB3tuSmKumPyAg0zBXfoxb+xp8weBQwjARibVlYpleh8OjLl4f6aJPJBCeP7/LDWNj7m3oZxAC
yhaQj6Tzsyt3OvAGDERP35GmEtKAgxYo1QvbW2wDOGw6A/mvSd82in0YmrsXXrrfsKIjNT6du/zI
xvu5nAZXqF8cNyeF52Shjs8XN2tIxhaxSUZR9PN2j3NcETHIR/F/X9VXrSpfv7GSDPApBexO5ECC
rdAhkETEGr3RS0FYwWKStKCmfzlPy+Ief+bMbK7irQbw1FrCKbwaDLE7rg6yN8FEzOSz2IRESebz
PY8z1AE9/pPvgPjA9a+Tdd/BsPFvD6D6lALZx14vK1hnlWH+tnGWuhElhcbPoni/JYCDyd3/gwwx
RLc4NdYlo6c+VMv/BGqz6se4qYgGSjWbW/rvkHolfpSiXO1cdHcj/HK7yG2Ksxz8MjfbclgkXP7Z
Tm/aD8MYJG0eRjSqDRlZiUcws9NpxONf5Q7HwFOu759XMyioIKzxIYonx+pMlQzdxpI/89DZx/I0
5uKe+r+AFZK4KJQ0UoYSOZExIRlDr/Qzfqq/+lvjVroe3MyOcVu9M2sl00LZcEKCLcLT4JDkh1UZ
B/oVeYTBPX6oSTbzVO8M0TvZNOsXkHl9Z5lOy4biJCLQQ3KZqeg4z/nmKLwWiZH/08y6fYcODpys
v1AToSKslQvQhiiASgKXmrIY7ambGCTKeiBrrbZk6DkqU61IOYgYSAg5+JiLX2NOH29nQpfABZ2b
wMjuylxreHDxYPGZNA3kwrZi0vXdcXb9inlnhrrM8eO+j2NjhkKZBFxS67FzcEIAS2/XyeaiH3Aw
1gyoP4N8ow0mRiMOkDVfykxOwUIQSu4YI8Q66bjCz/d616M+98PnG8yqR610TCa01EnQLmkCl25B
kM5xBfKYfq+adhQZnDXY7aOzpw73TaCqFA4sXTWtKj4Ns//grIvW5rVsH1n7cq6Yor5BbuhI8T0X
taq6NM4ZOajOfSM2n4P7qBDQROKuKcy3tfVROLyfbmlcpGaP11zSAHY5rIaCdXYjDoCj81YLsiHR
XPWYJOJDhTIF5hY3kuWt1g0r7wMbNaqv09hjY8Gjf4o3bKHoC0Gh0cMjOAdK3RoS70xJL3IFieTl
SuNMG7puDu2csW9pAfImGQ8Bvrn0+mAkQR7h8ktoT3T9+Z8z1H1s7iykEqjO4H8yUFU2rgn56vd9
jltuV37kUcfYsLoAHwqjK/RH1b0EurdSWdvg8Ll9HcjQ/gHVaIBonrsYmAD0GmpYC6lHSWT6Ihu4
3RHm0a0htkj4aS93f0u/FMI560BO5triLJQGAlkJ5JGPEx5eegyva58uJtc7ffZx0HAJc17m4q8B
RzZbYymK6wXFmjyMnPqJyTygHP44+NPiATS0CPGt1+u4jf4DDE8hHjPOCNXDakVbdmESJW209eQX
SbG3tK2JY0ZLHR78rcX3rDgtzvJctEHb/PQk3s0o5wSrzxgwfU2t90+IiHw5mt/x0hy9AM8oAJgW
9xL/ScN3xWBAQphccfOe7sHr/YMrRL0pNAteoQp8pZjf8yWVW4bjOgORG/+DuMJLVxzll+xVe7yn
95KNN92E8CIGiNKrQPBGx4+QP99AP3C3B5NV2hjmRFf8dOhAPpIU9xw4SBvW+Ifo0EpsuInMSh0t
Kl7vcTVvIeaTTTcRbh1JJDsHRZq9KUBzRx+WmGf8dZSB/IPKtMjjgYQF5nuVNg6WnW7XcCM5DSsA
grc5kJXAX2vh1hhCYJv/J/lTMBdWxzFrb+zsPZ/k7IOp69qkLzXpAkapYyiIJw+/sV4UyP8B3PKH
qBA2+Es2pu2s5cJT4sbgyjVIQxM8/Uohh6T0xq1bkVB0NHJ5rtAWEogGPfD6y9TFh1v8Mw7N7KPE
vRFhpxBZtX0QS/VmPXkVKAn87gJFFTAtVJbIB1Xd8u7YYUVI247dGMRkWklUJxn9wN2OVns/Dbm/
51jKY+moVM3uJ746CZRGWq8fwf9JJzDOZc8qdkSVre8HcfMNc80y4sU8EHcehef58fjUCUsNrCHe
PNRE+zrgz2VzTPn1oDZvR9KismcVoaeFtPZluuQ4pgctcsV+9krTtvlMF8K+pv29Q44Jlt/tLAu7
sv2EZTjaumvwXdGGQN2vRyURF6TURFemdUscznKAat6vi3VrpNZDH56kdw6GVUZmKg+j17j13oUt
APKyIsKhhk472NXgJx7yvod5VpOSC2qWQv7Fn35hY7k2zBrlY22WTNMffRL/96JPk1kpYycGhvhW
X0lcSAIB/1ThHTfwD+fm6uVfa6DREIdBdsbUOZ0Ow0H+GUcX2AecjNWR2z6oCBbadfTGS9B6z1Kf
YGLz4Kv6TnTPKuNE5G7WxiAnYs1Sl+Nf7GwSxngxel3vvB4aCidqOSJGD7VCV1OEWJuqb3iMBJS5
DtjV+xjHJRWbWl8v6ke4jRMHACUPewW1smVkjnAvLggc7+utw13rmnb6UtGv1AoHpTZtbWommzYt
5bNmDPt8SB9hnYZ3PAvimyOzLVFbu0ZaqVcZ3ZOAk9YB358MdFt6wz2fH4nijNGYqumxuBXI1IQG
kPdyT7rnwE02rPoh4NmdmLwuGZrVlEQF+7XSM14y/cvQGHErejLewydtcu1Id9cWnOH9iaHrWeIx
EaE7pUN7frQAOlOgzoyx2RQ1FpJtHYJU7gzh07oqXaD6u3ey9phXM7BVF1OMaFrmrPId7mvm14+B
2Mye7H2G74uV1GwV5d1+3fS5u3cNchXRxjO/S1+QCPfptSLWUbpMLy8I2WTHTiXQA00/raJMps+Y
AXfkrY6LRr0/saBf7dCizeqUBiJp5kigO0SvhA01LY8lS4X5DbWj/Th1TDoytl8hVV47w8+hc8wf
L/XstV+B9IZEx86x+IQvhJD+CjLFmuhvw5ns8y+vbah91NIQZ3zhDZ2KC46zQCGPSDRoZgDQ3XOo
IlEY8cXW/0uCmjlnT4va7Qa4j0lWNrUqbPhQhu3bWcGoE8TUvpgk1P3YzjQjY710Uj1FsbbvDBkU
XB1saUr2pWKxzaAZjhkCZwVCSYiCr6kxyuIHO7EPuMjsdNNWIqeALympG14k3BC1DTjAIOciUsy3
+6d2qJagYYXlNBItrWvm8+WBwSlJ6hFek7ftM7J/Y5iTcUi8Q7tN3fOPNcL04diq7wiY7SfMnM3b
Cw2FKQ9xr43W19FfZmZQ/pzZ5xd5tJeXbL1hyWcp4upKhjKuA/k99cVWwvuCEbaURrgb1RptQ4fk
2wf2y/x8e3qKSpWegkSr4aUuQemafT5D6W4NQJ994kybSMbPTyGUZ29qAPMLceF85dvLOfQPtuf2
yM+kwRP3w9Zh31GY3J0LebRD1bFTn5vb17GarSLvfygUdnF6bw9ZO3Iw+SP/39L7oJkzWdo7TWAm
MpYxJCSqwl1YlZlNELWcuOtcyzhXwXSXb2an2dovMc6hOdyeFpmrr36ohXkp0c/HehOYZwQq2kTN
0VGk2FoxcLnU5oEFOq/bjTkYF2fPFIYJXMpq8hrd6odyi96eE7npBte1nQyniUh1+uC8dMXQGsME
ShwC/8o++JZHZ0s6TFcyr8wV9rzZNOmsk0lPoWr/ydPpQ4Ilu2i4XSoaXyqGcuURjP5iazZst5Nw
XOGq5YhgSrxwgngPrycIprOf0vmqtwtVIeMGzZ3YgQpdM+QVYUsksRGVxkyo3vKgFqANXuJBGdhI
vgM446dp0MH8zsEaRlN/J+Fh8Z4uSkmeMVWFxjNm47X8uhSObF8+ePmF8K3T+BPbW67Gykoh5/CQ
OoYI/LxKXQgIJ2E82VnqUUcJP94DUEsOvHy4X3pkAwv0Ir6uo5+ldLhU27wLgVBIZBiGqPIZ/Yha
MBZeXVrWxpOZqJlMtabsUPdQ/riTDjI7WrfJQkY3kF99eceawXeMUI2i+JjDwSORsxe477qxeNPL
3/wSUPR1trOg9SL2wg0S1gDU2ErC3mGWelIVpC2lIQErDllzLIO/s3Lmo44uyHXpV5AerHlCLd7S
hOjP8y59BTS9U0FdE+DsXlqtBLqpYTdruxvmo2bLJx1df3GuB/pwiTWl7KzvYfD+FxDLW33fPEB0
xsRzBwyAd4yXeWw7d4HBiBg7f09LQ6BN86lTW41yPq5/zDf/w5fHxatVmTwZiFevqPAs8DHBXZPJ
bd4YrSZUWN810eeH0JmuxPk2TwQdcgIHFCezcBh6nex5ZFUezT6VawUoWSbPvEFELEH185mxsNJP
sNj17XTvUcwAjiyE/mwEOF/Hmd7AJFn4tvqasm3jm8iHqFCodvJsRTERJs6Tl83i6Oobl7e7APRL
6olZwKMmCio3mwlbsP9Mzgg84Ianmmh6Tz0aBxRNO9G7ilIB5uAfajm7bmfmhtiE/tQvpnRrbXhe
BOH8XzJUhd6RZ1J3WHI2hf5AuROJCck2PTBCP1/rS8eonQaciUFSFRPN041J6j2Y8BnUZJ844YzW
wisoevFoSjmNv7ztDIWpRYS+igXahBHrwCYutdqv3cqyNt9BxISHQv2X3TW+dIYODAj4lS0OSdOi
YGsd1DX+GxKt5/ZGZH5I7ubFH6F3pkMk/9Xt6Y86KPQ0y7yGHmQJuxxxFHjao7UYRo3xFBSPjuZB
FzyMm/aepjjYiMmcsAEy9ntgju60x1b2iQLWu32Q2/SdsDT0Z46FoPlVkkC5oizEQakWpSn/9I+x
xbfSkhTharlNnhOcYOUGZtkTMap+s40O7FIOeN7tJvQwJorMJGQKq8JpDPGPYqZEEvTbBCLi5MjW
ZIKOkO9yaqoiGpZzVoJuk7x06nV25JS1eV4kxG98LVmHRRuCb8idY08EXSFCdMGen3IPugkG+Uqs
mBJVXwSn/Kx6b+kgGYABkSMLhArqEbcnu3kpjmcWr8AcnjQC5fZbGbcrqAlq7jisQsGoGCgPBgh2
LlLusPYiCZUC2QAl6Js4MoCINpCzIET0xlFci004biLXtCjxPXUfG237044KwBOv1EebsTT5BZt9
7U13rLRUOCai8UOR9AYBpLaaaNIc8U8p5mWYuQiHKoWYMVMcn1/6S0nk0N+Fdo96yS4UrkwxDdFP
EyhS6NBvtC6uKdg78qL/cd9NoPCboCSjwVOFbGmPXTMMqF2B+Y/feec4E7q5Ycp5oBtdkC4JGnRS
EEscOZxzii8q0k8PTnnaKJ5yiKcNaUsvZ1mnLsEFYrYe3nvOiBK+jzChw6ROKx46WrD0ryxnVgNo
YRNzpEaLghWfw1VNMI31cvhysH/P9HkL4qxOWr2MM76l1rY9ba1XnuckyK+oF8Z6ZrxAMnixUefx
rWrP80PlDCoI+DC1AHGg65bBehbQM7SkLnt/0qyJ3Fn4mQ/ROfxgPwxkvLApUi8NqKGgBV28h0ne
TF5G76c36WnIzQOAaHMRBVIL4fjNOCqAP2gp5ZvH+iwe6mlAffxjUq8zqflg/J713ClELWogKJyp
v9GRiYoW6Lim58OXhaSzlLRvbiMFuCBBMakH1hlGUD7SvZ+5m7X4du5NZd+0lmw6n/PC97QbYej0
cClYn1iiGuEEZBy7KOV7rNtvxSgQaa8uc5Uhr69h76BV0Rg58cjmT9viTzNztLhmMzEhQN+qR432
laJRzVx/GU3EpCznCXu9eZfiRqV0hTNlZvMD0b1w5HnWmdagPq5Q3rei9CaYTpc37lG6ntPpzUsO
7kEKY3G3VYF4M6iCOOyq7aT04i3RFTh7U1Qrum5rsImmpP0tstImfrZvw8dNzt1wChT/EaXTKbEu
kce4aGGZYO7TAvJ/kGIb2xh3emZWAWm9uyDFdLbOktvTTAxmcgXc+M4NWRuPwjcNmarDY+hhN0oZ
2ljw6vyK5qojuznqR66w3l9+y0DigkUMdPa7fmZ/QlYZOS9IVZUTtE9DedmtEvpIdr1g3Ld0ymrv
eFU7OOCtAmgBwT5Yc8LTbEERPBbOLF4eKt5pykaZ8fm5RkqQpY7tmd8LZWD9KzhgEXnOKw8U3WCH
YHyH9YgDWl5fFg+zxbSVzeT0Kj00isZHbrpLWFN4k3NlJV1q6JBUKj+9vphJMXY8Bak3GoMqbSoe
Om/3uuOpwbzX7dYDdJbf8pxLpBLnG1feHWEdCm8P6BwwPS3a6mYHmFLzrevO6uLsnIHMVV5jTJJ3
uwFdJSYQ+Iw0CCar4rggMOMjaxrXTVD3IDVqraSpJ7Ws2tiEQFvLaqKm1clVnS9W0dSN4wWvAcIS
LczoPwTPXOSCXZ0t/Rxhfq5J5mEk/NYO1/W/G+UxDZPf/6n9r5ua/eVzk/egsHCTz7VJVuQX8sWz
SnUmz6RkEMrQDTOkmpUwf+CeylZ4lvybxvx+NE18b+DCKcLeBG1cKTZUaiFkaKE38U+W+mR2j34E
82l4JMPfHP+/UaiPKYNDYT0ZzsBrFwbwFN5wNx3rFYS4S43VCcMb/cOpAFPikR4KOg5JWM69ec/S
OglACj745pNSO0Qr8UvlI+AKx4fJ7ycaW7kRl6HemQeGV0losKtvhhMiQQP3kZprgPJmZx0kQwcJ
+CVYPVxfatiBYaI+wwHKzQvgKwaeMqionExRXg5z5TI7Sj4lw26vgSHPNnGiHomrRMzpDKF5fPvV
CRe3QSCmtfUxobqAOnuM5RvCEB6Cm6/6C3FwWFgh6WHA9Ea2jWOyq8JB+H/89WbsriCJHSiZmHbf
C+Hob917aRXYf7AMcu/xtcA0OQmoKxYyl7TV7qL1OKt3/JoLRLi0DBB5wiAhp8p6GxgUOLWS398g
O9+YriYc4kcDzu3Qwsuvhq6QuYCRj3K+Tzu9m088jUIO8WcupHm3nTkUz7lIul3YwBHKWPFha6cZ
Y0EVCbIk2CYlHp6MfEgC6XPWD6510a1+bbo9Q8yHAIkkAgRp3h480JbeZWNQJ2cQY4sh9SGVV5oY
g0nIF3k5BxLvpKansnjGOMJSGCBIOl5pPn8sOxYjF8criebUozJ5kmTZEwmnQipELhNVXobOapIy
Ov+P5eXSy1bzwUhKppyrtO49dyjSzUzbabwBRun4Q2BFJlW4iB9iy0QWvMWhBVI30SRgFPN1pUym
K56bFQJjJuNv09aqGoMGx8yRVqqKRX5w1J/9A6CUsGwaismH4nxxkf2XWG1MgD95QatFnyzkHp7J
+o93duS0CpdedzAxuLgqXZm8fLFU5Eik3QffK3TVCSncnWINuwxBho2YpMSmzsrF5cQrrKis6fmE
pUJSI6K4tT4IhLI9aDmBcL6omHA7aJ4Pbz61if/S42aTo/j7+uyAsrsWKha/Qd7J5nEjrLOfQMoM
gZdFfg634bIDWv2nG3jcX1IELz6pTCt5dEyiNZNdTOqZpl5YKV3mHz4QAM/2gqGxqJ5qo14sWa1n
CvWvJtuja6um+iZMEUObtpH281x62ybac+rXA1KjI1HcKian6SxH+SvJnD9hlvHNTBCVVuia6/7X
omBkmO4OdrLEDgfTtxIrOaZDvuichgI05vDR1sR4RHknGI6g5vTRaampf4sa+YPkZRC6YV4cSV6y
2EsVxA72jnY9PWI6Dfk7yY75Nm5cphEmqBFkVAv/m1bfPPayYAE1njGJ8Yijx9LzGvFVHQEy0Yt9
DXbk1GHY3oPckER5jVJmO5oOgIF8SN6MkbWJopQdm7haS9ma+Yyr64S4G9ZFYybJeZ8Odwc7XjBA
s2mD0bF0efw2QP7xUq1s5eezWNSVV0NUs3BeZ+qlR7kLAHn+hXbGFlNG+5wQttwh2mUnw83IrvDf
ThaOgy73lY7TAdxwCMK/Js3Epf/BQnIxkp7hZbqUG7K0bqeuIY1HoZVS1PQGbf17HMJIoCzo5q20
3asjuoyjSgrJGGDobh17leieZZdnlkFO+D8E+T4yWekAPSvuuHau1/fWaCpXxmT1uc9MfSLojAth
V+LKX0YHUGsnD5Pm0OEsHuK0UFFEO93nXl1jbn+GrbWz8U89qt++bnp87KSsOTNcaAoJnCb6HCbn
crIc40fkufNIr61a86qQJqbinpyDt3lhlWNxtqmgTE1x6CICvN3jTc2YInQnsmpFqjFvixRf8uc0
uI8Gy7dWfN6NljybRoz20GkG8NI8aLv6X1qiRtpoRjdyL1I2NcDGR9/PL1T9IQsZgj2/5OVmFjiB
PK+iiVfe02cc+beSlHrt/xYd8RXzOtZ3lX2x2s+SdOPR7BDD++m3K1CdQCoy7Sdy5/3bwfv7DQCS
RHcmnnGDifRGW1J4zWqfTBj91Ioy+TbVByrPfAi2ADRMTYeSgkkiBE0wtWcuNIL+mwckGrknhNjK
9HAyDL5/gN/AtETuDxccGyJgfyr8EmTmdWFPRwmLsZW4DdzkFbs+6brsOfVC6UbmoOX/ZcluGXeA
lUt59bdF3yg/+jbYNVxJcxA4CaPoFEH2s5DjNH/zEALEg/A4K+M/vqHN0NDFgioK/3xXHggPqGYL
zAiaElkWxG8CY58tnN62c7ksSGe3oIZoNLcOWWW6QVFQntdG4rus/HD7wQKloJgOR0jvYNdej5l2
QJG5iMKv10teOXKVGo16gW8ueADTMHYZjKcxORdgr0SnkgqzVnRDzueypzJd85iogGhzZ6MqD55c
usVnZQ3tELptT/Nl4gWNh3q8FiO4ac8WM9ss6dNHAvgASBWyRJtkZyrrsP3HXGxTySFmDlji+pIA
2ceOVzEcb33OmV+PP1XqNzdxn+uY/OdKWEWR13bEWRntmGZvTTw+eySUxhROjp2pe/arEjOCbfTY
A4Sm74+pBrjxRstx96oClUDoTLT9VNy3vgWtpCosmkFv/cqV0KWUqMxCGrdBLZl4AbdNZIvNwoJK
ZvmvweCettMlJ7MCH1oxRDdrcD7yYphy/BWemp1+xfV+BqgqMCitL8AX8GnOjMzDRDZ+fvwjuzAE
R0sHCqyvYTl+4GGjXENQFAImw3oP02m9lIWfYWAwNBlzbknCD80g373R6PxZHlxP53eOcRloIftl
zd5ad40HPipFiixVJp0PI5zpsxScKRvbJu+pmovmAbSvjOt9nR9gxCVy7Ryh6FpH0J9ApU4pZ1kS
neHB6mDy+4+3a4AnyXba1ApsFnuVMcOuk6MNIQ/0zKf9wcbiGMgvOVC+jV9F4oEUS2A5s3PZyrpa
y8YIh+aq1ceWhWXAtrCIRniqG/ljJPv9fJeqKJuR7Zlx1mSb7fPXdQOiykw9IUQmmviofbDA2POR
XLkkZik2vFJrHTcXYSEkOIlQfruIqDT+EfI0HopTHDdyiHAVBX55hlj57Jv85EyUiGBQP40+UlkB
9XE3/SwNIGF0LMjBoHK6adJZ4Wg0vbl4rbzHs0DB34q7Bsjq4s6/6ERe79GqLKZQJ5niil5priQ/
Bw/x0KiT7j3wkCBmi4IjcigEMRgURzv8mD/PmdpYfg8pIgsG++tyIGDhShcMKxaG/7qwX9CaYiEo
vU4L50BGBwtd4cHGYajjMgYG7xfZr7nNikl8SmbjpsXpZDEOsf+6Y9TPmgLgm6ZvOuHZDg13hCy9
0zI3ASVEY9s79ha3dC7M5h3OCfXDur8jq+fyRmlgUNcZQC+o2QeaDwRAUkNxnrxOcaEsKgssmZKv
5er1ng4e386KLvbvcQUfNIkRX4AVHdzOdBLer57zlPZ/a+MSx95UexCixabxAEakctO6VKAyq7Sl
0vh3A9cdy+pGUdA1qnxhdM6UDNlVnaMz633n/AnIqtpdNbMnW2OAAG97dtkASkFGU9jPVOgFkHnk
G6Bb8SxSBt5/Tcc5+WRQTqSCu2B1wm/KQzdnOC086+rxBamd4FyZzgpaw1hWu+cPq6uJnt50WmYA
O2TEIonPUSAP/3KhOB7aczKmFDD/rTLkZWh0Ddq+uaxaRIgub8rYOkcqB8bsh7Wy4MGeqNqv7m6f
X2dOyIoZY2tWDyYFso/3bkO+3gS1xXWzhYDeODI8Uv1+QgJ4EYMo+q26uG/eGknOAP05WTlE2MfQ
mUOwuf6gplfbWaOWMpn8rEJ6AVujy+KwtlCQDk82eMpUx8u2+fCzy2Kk++YbtNevQTv1eKVB0+Vu
fg8d2jV/BtsrkUMx49Ie897rdfC/mYyKLbBoO/0PeMlgbTmpAmII2Wd7RH1GiJlrVPplsKh8rr0v
MR2LF/O3p3mKzn1Go49bKiXOxXTcJeteKfo1qJBI8/9m/jcWw7IFLE91XCj0+gq8mgLawDtmLSnt
a6f3pv+Z9bqhGKmsUAaFQlB3T7jZtfAtAu2mzYb5YpuUSJ8PqtHUS8PjtbqytT6RfKDTiHEwiIPm
8HDtL02VXgYfMYUye7iEKxeUwYFkpp1U4uLx3HFY6zp4gyPTjqBYbQNyVA8/45hcIQ5HcLAb0TPf
LWpQ9X7xkMStNPiRZNBOIB4DnndQGsE4ktiQS6cBK4jjdT9uvyzWabjm1ItHF66OVsMIKPLg1J6Y
LU1RMm7QEvbQELzSoEtYwR6b+r25IUjR2DBqRzuyDQuVAkV+cl+am9bQjcsV688bTDommzVomayz
Mg0YvILFUxJ0ncSnLvSK7fxuo/dmxzkECQrHDaLYZ+zNyJaxMqCKKAwdahVrg8R+qBr15j9cn1we
SNq+Pq9eHhFemE4NPzAyawJpcPYVAiUDM60kPppKIDr0bB/DYI0rjD1tr+MiAt5UPFLF/7rdMk60
2RAGZuHeAzkQehvx+I0D+AhJI13JCbEClbIhNAysF0ODxWUxq31ctNxgOwuDuxCLOx3fpl1purOK
q9Qo4oeUfB/pr2TO903V4zKIomJ8PUs1TDsdyKI4McNiTqaqoFjc88l1SzsiiJfvEbQA7Xws4uzI
GsLBOR/Z6UXtWdRne1lXqWGUtTfYWlX9YhXyIu9iX4AkrKvv0jFRKl9MR9uN1pYLpTmnf/cR9QP0
nc8eO2vHIISpy7W8ZZMrZMwoSyuSLhogUu6pF3WkF/LNvzaiw7xDu4iTp02F8q0OAhiNiw0U50yZ
xMNQOhKdsnZSwHsAbV3HOCBIvEZF3rU/WY3M0EH+z2Y3EQlkhALPC2UCmmmnZs/qqQI2+S6p1sD1
BF1gET5ys7a65ZjGO5CY5i6Cq/j50aj3JmiG9hjuHaE0FP0dfSmOAWbhVsU4s536VulSa7rJi/5x
wy2yfkQBs4hKOJht4RFzk6ux+c4JELqu2+QFvpMMEbqcumKd/9Y7jQIBjIJsBjmLCMlCypXeudHC
RKCDW+2DM6TrAtDe7VSfY+IKw0/H103zzA7eH8LpOMfarEOeCE0H6UqvdctFenc2Bw70+ZAD+Oz6
E66vXyDCEyAtK6DngEmk7E2oZTWFaKiLYDeg/HC9qZf8O6ekPxbRElslfRfinyo/T0Qj+o/LCWNs
kIraIyJDkbTs2tImK4ORzkhrlzcXkj5HLEkuUgshlZ36R6nlo5BzzfbgNU4tBGBdf0egKDOWBrbe
C3bzXn5rGiTNO6886Q4hBeSRigee0MwYBFqUU4BhEmxQHmlkUtLT0DxtvGeBXlf4ruwXE7Rf8M52
5yPdAb0yqAmD612GZoBeh74cFyAOYpKO1X+PcWLvnIRgRGg9MAUjeDDyA0h1KL1xlRG4HW8iUQTz
QZBDoL+cnmjD/CwtSZ62B9EZxaRt+CjJknglV+bFxIRPUse+Ds/V5zH849mwq0yzIu38x29amove
CgzwWLszZPmqADyWH0H/25YCctEfd8g+Op+jnVfDPji17CCwWhdx6d+Cl+FvlEbMUcIVaP3aBf/Y
7D/QqUH5Y3Uzljvb/PRhPYKsbsDhyicP8o6k9AOkMIvoB8tpAxOrS1EBiMFY9wk24pF12eFhNaj/
fqsdSwUD4oMmVo10EsxT1vfr3G2mEt8CwgMvsod+LKJRfjI5puXhKZ/TD38L1ORZbbMiu0MvcMHF
7ZjU7YUbPB4M5Vl0KE1eSf2JHFTrvhqIIpENIlEpgM2BhCUiGb0pDUAV3F4xQ8fXYIhnnRU+Q3Al
4tWIMVKg+rAyJzFbgGiWP/9YfR1qFGXn8M4vY9mWRNImNPZFTUWb+vm34h1S+vjZCBA3Cadu7f2R
M2YwAMeQKZniOowQj9mGfBNVxO87zqwlRfwK6sBWYbAYE9vBTyLk55D+DQx1zUr9838D1ejyfPDw
PBdLuTllq/btqNibJ0HGQzObPaNoaKJhW2VB7fmTpSfKIokILvEzpyjZ76+GNn+Usn+RAVZ+ZNTI
hZqb/T2IyqJVYyQ5/pSS75K5m/ucUZVRdMG2yMXDR4omE7RkshPcO4pPY0jbg1YQm0Y5zUpppfMt
Mo2eTYhmVr6EV+KNp7A+b1Pgm/r5nBykbs0Tg4klzNlGqi0maGilPtWxjClW7NYfpVL7T6O8e/Ru
QPyb4cDbYnP91npZ501O6SnmP7ZFbfTUTCPKVVihMMWYpRmh8bYKe+ZxgMVgVQ0MR8k8tt14Tu6Z
9PnucIruyq8e3O1MAWNkto9G/BtzS7TS0o4mXB5yNxlKb3XY9RAh+7QK/YuiTV0x5+IAmV4jGddz
kS34eiJ2c46GhcCLnKP7GcJ+lWRXqS4IOn0fFi5ncdA4WWxI33GVw1wLvxb35L8V6o4ubHIO5M17
SBDcVauKMHZ2BV/Sw+gopG8012YF76WkVQyiP7F6FqLF0PxEQuQMRp2KjWWSUL5JjCn0e19SQKd0
Kz1+3lyN6HgibqX4n9eLoXw4a5NSQPpdCxFsAFXFcVD3r1iMamHSU9/J7HvWH37mcE2CNS1kyoQG
CKaXooHetMN6bjtyAIV2T5K3Ei9Syro8GY93MZa1TBNSOx4bDMXly6zE4pEBRKKy0JKxstKNBzss
tcpL5jKcoeFZhGWlJoyd6i0W0QFaqFbUZa8JY+NDXK+egipC6JhSiwMDB3cuLj4jsyEKoQGdN54i
0IT244BI0hDQVlV/zLSCHchTNuvpgjYBr2IdrCY/jsjyjhmCXk9RQ4Jteh2abD7oLzpQ/3Dv39No
qX4glbciv744/UTgdbU+o1JXPkQ0fZhXHrSnaRmdXtSjPbGlQbCAIPMuzRd4jZuFqUWvkf4Mjs3P
48MlgK2IeMYDpYLgwF1C35414eh+eKDsS4/YmDxYLPDQMoXS74rxtEK+tG2SVoTvEdkz/WEQJQOG
uXtHGOFjDte0PzE0wCACFW8q8igQ0/m5kOULVEwlqiFM1m+MZzP+ml4x1qDLvqRZHGFgToP21uYb
Y7RSd0177lLWRi/fu747RwXiBiW4NyNp2nbOU4Sf8SBHTVYeDfDU3Okva1n2X4x34p2A3ODBxdjQ
r2haSeRW5G4jDmSkfSBqujz2lc1RjPwNKU+EG8aGNTCJx/np8j9MrjWN4e/A8BCaxNPSWWLZ3LeW
IDz1lqfG5GbyqsxNOqqm6U0Zr0Q7oks+t63SdOcCZznnHCxxskfxBg2uDC4wLSn3pAKHCwDY+DGW
ZN7jgQRpOaBKMg150J3o0aKzUvjMiH7mgDPHqbByL2nmdr7TolhfC33OODihfEYqnVarG8NfiWGf
BdtvuUxd5vBvmJHe6tYRuxcYsXroVg76k7XxVwqb2t6r2uUcipx29qTWPGSuhTQeUMoVP09HKGGm
EWCm/XpFVBdJ05u7dgyycNWkW/mnHF+8ZZS6euLZZX7TE56o9g7zTtASv7u/W3yex+xkDB5VDLFM
0jl4RoexdE/k/gMfYGp6g7MN0TL3acm4baLcElSpxWpoCNfEQbn/W09F5v6qWNvmGQjt989bcn+S
USk+RrD+TMzuUqBoLuCB+Xh8MVisUG40TxzMIL1hcC9wsiwi5MtSi4Dtv9yqZuq9rZc0zcWZmr89
bjc+W1fxvxKZCh2agFq/uTjwI8nOuxYSIemjD8FFgNRevknP/GVgM3O3DBjYq2IUpkORemykm7k6
3+pJdr/1y8pfsfJ/+TZV+2gAAtaQKgAQpj5+N5kNtCfKxR03d0f0reh/llnjyLsvmy39Zgo+OnYc
8nXpXsTNQNNrxY7DR/FcQPBBnO9Eq0iBbZ6j2Y0d5Kfs7fCaErxTwsutR3tOB2Wljb1KMpl1hUog
mZkHul6kDjTEWxWxAa7/cT3jkW+3c+kXWCNxfVX06kKHeX2KabAP0v85FKKVSQD/EG+irjQwREGV
N/4ocOZL1gBb2fKozoRrq4T3GMRvT2mY6aY8f/ivgZ49Fzl0vLTLHMem3VmX+4hFACzBx1+7GcxD
oOmIxs6enT61aXStq87V+oZt9ing7tc5c9KqkgZaNu1+izw57spfBRRCIgTBI+feWVgk2OuRd3mA
lkBm/kUpGIWFz3iv/8/3mgAQB17TEbg7ueOR01Qj4Jh6uW9+2ho45lMIrtUUwLF8dXIQdub+ZBB+
ke3wU8pBHX4IrGDuXz4xjQTj4eMmsibOU6bppgxgoK7LNHQW63vihyrU7EVxT9ftowCkSyb772Jj
cQnPnr6kQC2eBaTcbicOhwRkb7UJ7R8PUQ3guo/dos1kE/bLizIyQKMjO1EmvEqeDu47hVXvPd0n
En+DYEyScPQ8xdRksfRvOr9b9nvCyvEtUsh0oPSM5fTHfmqHhYhuFPa/rTd5GJ1ZzuiEWp0iTEFk
6CVOJvijF85n/H96wqEP6NnjGhqe6JA4R3/BaZrR4km3JpsmvFyVFnnT/TZyQ7dxnG7DnjGdPUJq
+NDlbv9gteijwWx+9x0/M+X2OCydo59LgsgyzwJMGSx0sPl65KgWDzT6T8UcaxItdf4n5UEs3YcZ
ZNg0or81yixkzuznrseHCIQF75d90N/eQcGjZGed+PCDez7eeiNvtMslivKpLsRil3vvgo5PNzyY
TftdrC6NpRzctAutKJX3jpHaMiFUsDfByg9f3l+liYmcuB5Cc5OcgSwNa7TJE98zKAGPR+zgLi0q
TKQmYmwwfc8/giVrQTgRERPRbOXP7ZVlcJ6ZG6MMbfOGqYnC/+NjQik1fpclMO9w2R4wevoZCNt0
eHq1Faz0HP+3NkP5RZmsw73zUPMMKPTiw5cNY5rD+nHSrXsjLY9xirstXo9eqpg+4zGCbw872L+x
irf8qGeGqwdYP20EdHYSdwuTivMbMInhKhhJcdzH2orA0JYbFvX4HBpg7DDlYMNJ++LQkgaDR71u
b82dFvGtTOVpDXX58DTrZGY3dcYy50l6moSMLIBIC+OZ5L7ZVj+EyAMPuoCazVQNB1a2eHDckxXW
9dzYB6gqAi9DxWJwoY/tw6qn1ef1QCdGYF9esxGZHgSuAMYf4O7L5xa4dwncTt656inDW+D58ajc
C8m/8b8ocHBQu87fzZOncoS8PueLQfj+QZiZRdL6GH/krH6+ILpkg8glRDYuIY3+07/YJNmQdHPJ
2UkjfIoFrQPCrq9yuCTKQLt0TwhqtbAG5ANAWKFisvupi9PIdMCqt9IdJMM6memoIvzmZ005hbyg
pDQkIYOM++RLhSr9q7kMCrciT/JloSZQxxkQBOaO20j/1i/62HFgnlPAQzFsXmoBRW1dSqRl+PPP
bBpjkosDYu7ZANP4dTGAExTkcPxHEh5TMloNW3849NAScuJb7S+szaz6f7MdtiuniJV0QoFewubO
HFwsT5AnIrCD3PjDPY7PzPQM7F0m8H+0oARYmadoJbyfcrbp2+XlC+zEAH+tFCsAlq8vsV3B+9xA
rwOQckCyn+VxLjr1WWMvO2tAurMkJDmUmd91U5UxOJdZqVF7r1Lt6JE+drFrIzT1zuUk2/18AP3a
HY1pewwjzZkBShSI42UqrytRM+2VpdkqDJi/citSZ+2codS9Ftku7lK+v3s57bkumihpqFM+5ykh
qqZbnrSpaP92dwn9p3gOpVJXbmVx6KBwwC9H6fpPWsIbH0si3b02FPhbOsIxHo64uokeUBUeu6vW
XiZbDaLXQOCYwjb4ifDYuUqs3bhSE7zRkXxcOjwP3ERamqlZ9xURwjSJLZR6Qs92FeQkGuo59vWJ
fsMCa88iwk8vGCYUXwuVSZH+YHezwAUiR0mG7YwxBnAWVSAvzJ/j+IxgtjJRbl867QJcnX0z1g6R
b0BTHJa7o9EqrmhSvhE2S1isI8gsaP681f4VSBJsKJ+qLWFxD3dUNxTchPyFI/MtIQ7uRi7e45Yu
BW+t4wehL9lYeWt5479w3HsMkF6RJDqQdJvP881fcEyWkp9vwFjXY9X9eoD1jttO8uepFITQKA/y
/0tWlxLQnWK2ScTwd6cjVcrgOQ8gj6AVyUAR3Rl++mA6FhPZQo1tBR/IAjlErm6OOAEj7YQXcbIE
w8pErW9JEulFwFQrrAXiPb7hS9NylaHkLlrAV96HsCwzb6A3blw3dHkspFL5MoneVLFLAAMMvrua
eA93DAfiGa4aM6WCTVph7seH0iDF9HtGgS8DDCtUHoP9T7ZJki8/SNY9VD6YpXu5LLt3zjmEVufR
iOC1sM+I1jTiZuAWUE54p0FcsUaNnicPY9vLVre3s09J2PwSYScVQNjluH1OW768agYFJoGYlxzO
454EN6Z38du9SyNoiiI6M8aPJtsDRa0hlA/B2jUY+7kKLo7q8AWD+hEkhHtCFrxp5AxuXgVkkAF2
tARhlyTFt+T4PlveAaAuLm06YCboIBr8X3IbmGA1kFWw0ti0eXJbH7TqpmOnclV9cCPDNZ+iTwf8
5dveUyh6J9pNBvBbW/AUDwW/8Yt7I6z0f9xAJhQzHi+BYfkNUiF0pWSIsPCZZGdvD7X0M9jV93ry
hJLw5ojqPommzmFcby2XFsPPWKSmvLTY9CM0iCQSsQDdMMWz+3uPgAqao8C2tIcfnxGL8nwNxSbB
126zyCUyfvP4Sqp+t87RdQz10W/E9gs0JbLfpCJ/R2aqnfAvmRMEu0lutBuQLHcX0P3vG4RLj8Kk
S0as5Jz6H0Q24R71ZHUiJNYDOrvtd+hoZ53/X994j6tn1nNkowayJtmfdKgNeODiDRKIt/cvmNbJ
BBml6+jhCK/V8UosPW6QIs7E+W8ieTMKiN1nmbAfJmXxzWL+wmvv7njgESJMrlWT8MinnOopLkaO
Ri/B6oOnXKeWXUdU8yxjIAd0FXXPuvQ9cJDIwAl+yVxoUAjVYAdSa7CmusbV+0VbCtddntHNXBby
qqKJwMEp3hZbqx0Sj2ni5ho+/UepJGWTYAQgqyofI1G+w4DLvu90ifdkEzuZ6q5j6MeIzUJffEvD
yMWIK13RQKJm1lvtZGJOF8/+TFigsg01x3IyEJiGBgE40zP1SQBEpHc7ngAwGDfD0jThkqz2BWD4
oQmPm0tMW8kpzONMuVHXciMNpVYNus6bGIeiPKpaP2sXrN+gruepPmSHeUqSDfVhSQ7mFnls1hXT
NqLs/b5APo+EXdKl7N33rKqEZypUqWPjcOBk0XPFerj4NOnhEyZRPa8PwvVmyYLB3P2HfNQm37EK
Ot4TzrYUA8Tj4gHxSdTwfXd2jw+WYdQTC2G8kGNn3mwadOG0bvLBKFJLdU6bhcK7+iI/8XoejykZ
UAlbXDN3lEQbE65trCGZAEpbD0/syl0tEeJUPL4kbFq5fQQBXia53QSPc9Kt/HIV2Wy2VRcppWHS
pL6p+U+6G/u660FuB3fY9SezMI60O0mweydeqEojK3BRw6WscMTRI2TgHLOEWvn/Jfuz2q87YrJy
vIUQfEyiGLj9AW+cGvq/sQkE0vLZnV46BJDzScfKxMnk28LT1vfCyQyFFpVpH012xYau1OiOZAkj
tLvGaGVX4/G9P8yROBnm7P+XbpPvcXHpyyGFzgAX8Jd9lMytaG6b7ZioAN1GrxA5ORmUG/wkzH4U
n2JHw+7FZP44YnleedXMBP33NSYgFRK4lmmV5BjI1RxKkGSuK6je5MIyabYmSZodYguRboBeaXib
HqJY6HpS/K3uLr3Xej8mIbrFHzaGiXXihKM2v327ICW9Ig4X44W2WjSwyebUpmyruj8dwIF48cAj
ERmSReH73f//9z1zQhh2wTnFdEGvXrd9L3PEG6CNKtvKMeYoJL47hxUorLIwVEeMN8ImEU8drdiY
VTprS+9IFiZ/Wu04M0d5kWQeSLXOjE0dDFPDI5mgBAMQoGQo4sC+ApitLWEX+AceEuGdHcIX+Hh/
ks7Sskz4Oih5HvbLZ3VY/W6ZyhRYzpq9GsaPkI/3zVrAunkQv90wGwz/VMju+bdHrD0MB0fxZIOL
VHfx48J80soJrfKdwkD+6YeQd9p7FL4H2clREzm/6SQ2QmqS2SLqAmSbNnZBsd0UpSmb2b7diTtO
o4rQB6DJYqmaeG6JkCXkCOIOk8lX794xZ8EGJotS0OQ7gcd2MqNVebH6eUzhlQvZpTo7Ip+8oIe9
Q2apT1S71Ysz/1oYFwg1FwpmxsVA8VlRO1dJGJ0UzrRCeQUlwXAeFtu/y3bnx2/D9xgoKgdZlfto
QX91TCvTBsZt8F6tMiVeDxy9cuH33OR4w4p9X2LMd9Ulu3MgCHkg5hWtO16iMYGz64SMSxYWe3BB
R3TV1zeqYlP0Ha/mlJVytjELkzuS42OxAskaTxp2Jwez3qErAyLTEmbcsBvqXInOymu/rIpoKdaV
BKebGytKlMIaU1md5JwtozxBB5dVN5JV5/t3noeNHM5mKHdtVBYW+odqlrQhYiXuNx7Tt3hu1Adf
NEBb6Kw7G+K+RONiy38pGfz0oz05lEqPVqAhRjbulA6Ii16BqcmzT3dUIxnU8J/26EiaVnB1Pung
yFDRXM8hriA1Rys0tZnCsZye73VSYg//pA8JStb1/1nMoE+M+f2UwwzeikBQeimbmSYg/8fZt2Eo
0yrk+Z558F5XZ3bmCIz6GTbCWRopMiXquXV4VWf5zORx+iFh0WcpdprppWdBKnoEL/2+zJvrGLoX
TMFHMt1uIqj1NhhIVMbRx3Bp5dR9vpMmFWs84c2e3xkOeINrz38DK5gX2XOWh6evWnOrKUZ3Fszv
XiZG8Hbu5GiOvRYxFcylhnS+9fyiYrZlKW10F/Vdcn7pmfBS8+UpQ21AKDsTPAehOrkks2hGavAZ
qCGZxm0ztiOeecf07DM5T9YjzI1+IIzFSyESE6PBtvfM89i4DudOpSeOFeQSk6FKV4og+j6yH1XF
z0VW5mOck7qwX66tOl0LXXuMUI+hMG38TtAU5mgTIhVyWOb1XntNFefoEjjKjtVdaoaRpygWjD6+
aTcb5RIpG7Q3CJpgHRpxIS2QLCdUToI4HGp9c7ljMTNTu68EVcuPAUgArqlyyNSeBLKzqt0YyyVi
gK35oDDIJsm4RnuLIbiXCjVfthsye/bcQ3iSl+f+cEsL2Bf3Ji7AW7Qd66WOSSt5a7e1rIqvX6d3
uit7m1po1yH1XJMrQDX/TsYR4x4CXiJQ9oXoPEwKb2piSOTuObCoL4gYVz1SzddE27xCwQLCz6Ex
Yl9rIMleAQVucfrfetIlEO04li4sJzOAttzlghR/Oj2Y0JAZN0sEVKGrl5Cwedw5I9gTM6qxMamg
CY7VVYDenXa8EG5Ml44Bc8yYXWmrkH6taxO82Z6wyPDGS3ma3/3VgZNAWFxMcu/CLiyQXNyzpqz4
UdNkTBe68zS1LsWQI8VbPeDBIhRpgB5GoNtR2BzkMsXetmY/LEgDgDJH+8p7/ZYNMbL93R1fAW/j
OhiLWSue2au5smWE6DHcsvk9mipyeCcjuNFEjnGnDWjbKlfFiv+DDMLqTpV9xwRSHwZwAZXW7t8/
uUXAcTYR4/RCwtgw8ZNnJWa1Hp+geGghYsP0X9ybaqEmGCZWJXEWvg1XV9KIZAChm/Igubz53rHl
mPm1qhX7F9E9gJeIVIrzdxTG2GvK7u+rIhpFsXsSF97zrVmq2iZpKab6Ltd/ZPxzx/MxKMJFSbRO
S0qHPeLRIUursclTq+0vCH1nHXLX0sj7s8jsIf+TPyH2LB+Aap97ISI//QOzzNt2ZVioqQ4ETBH8
tOAW38vX0BSz6WMd+lAi60axl8VeLJekrPzL3qpeJaj1m4qIZrE/xpLN5Ck7VDCJXp36hSwIRidl
HUpcHncJt6rElq7Tkf9dssfmhjedmzjqe4Ow9zeTMkuOA6R8nNFqt9ygSzEkheodwgsP5l0ICM2l
YMQlqiTGBAezEe8RjK/CA9ct2LgMOQBHdHhRdUC+DYNE5c30sDWwr47zhQE/Vz5FwQy7uNescOyM
fa4hoTJcMH9lPT0RkztDkQDWrgrwzBAA4OjRajB8NBqed09o68P6pvWnfzbVBvZq2YREWCMwUEdm
x42gqTY36YnHOYJmWbEPtX1Sn47vQcK2lNOx3onz50ZcQmATDULH+lcDE4aFr4AdqEGDXE150yen
JU9fkRWtiQCUPMnCvM8Phl8vblKkhce8XgD/GzIqnWGBccV95AUaT8dSBi9idEv6V8Y7KQQaSQeF
w7KxXTnHwUxAIKqwuySiD8p4F2VsDvhdcadMrxSWqYh5GJBS8TenthJti8QFPSQgnSzNvzP1wfTq
3a6CADiOTOAH/loiWUnRHmRlLRJ2CMg9HVHBggTHg/AHuQlESgDJZqfoafMDIFZ6itOOYW/ADgoJ
ho60USLlhRr5EbMipvrs2ovHf8Aa9IKVBF/VNVhIdH5DCf2Aux19PUSiRHw30speN4f9/UBOqSX5
U08RUnb9Z2Oe221P9y0e3ScmGAY72RN6yaN5IMQmYPRJy/ZTHzwOaa7OwkM2g1RTS+ICu1POI6QS
t02lfEzP3JAGIg/HNuiFLNgIJwyBVvEBneIn0AfBT7Cwae0bOGFKlb3qtrmR66Rc0GW1iOsdbaIZ
Rvasww2zxfIa98jaby98rwNEy67wgniokpKxqdf4hx2RHBiLsCY5wf3zctfg2eUhdtOyTepPTddK
3sI6jYOlexvlXzhqLFGo5qVo1JQC9pAd32359oxUblyHn1H3ikmGpxLnj6DoFM6XZARmlCbjINBs
wYD1/R9rrPg3nBD4CQHHLdPtgsmLvyB65dGWn9+lO4KWptkw71sIHQqAUVYlKWE+S9r18lwZkHnL
j0t0LaO1xaQjFh5MrZDq/n6XFV9Dt+tQNkOKxvRC9IP1ViJGCWHvg5KstMHaEKxWTVJFuKOZ9LQP
JcXa2fwn13JMsdRkzViLWunIS0daZVswhxLC1lThGbZRWziUprDc1H03M7nPtpcVAXAzHpOkGb2I
q8j66NpSvCDbYVEsu9TJQ8dTO8MV/Ob5ETexsPtfRIszWNE+dHhUvI4VxoZxoUteS64RCTBvMvG6
HVKgMYMcxBQwoqkoPGTLb9N7OEoZGbxkn2kKai51dIIsihrz1lFodjjgAlwETf1tYfrEVxf/BVrr
02MQvMKcjJs307/q5TYO5X/F+S2cnk84TDbGakEtXRGHBJYJI2n8qODPmdSjNof1WfAB1OkjJECS
SwEiAn8Ph8vU/6wsYAslVW/YOvAddGI+x2buL520EYTPbneGI33olvCjxghdCcTfCDWUvvy2//ud
ZAWe4I2AoNYeiNn2xVp0zPdZEfZFYY9T0PZZaM9n7QRceAQW5uY1/UOQ7I4v5lLFuuzPjvI/2Ti/
RXZcPxThSlh7L94aLkhE1dA7q7ICJbTfE5Rbry2YW2hpGO5lzYx8tuTS8PbocJuElj1WBJbxAjcH
Idyi3t8DMdxI9NUHKFRNrVgiuNHG0v+JFYCrx8wXBm1UiQDD7sEaKDN2fXdgpSOX5eHxS9JFGmtJ
602yQ41v0RCxM7jTA0BJKkpm93wRuyCO/HcqlZ8RBVwgiEDb0BWkayrT/JpQ7Ob9XiDrI+7kji9d
N6ImvJBS1hK7yEhwKve2YXdIAbqgq5Z/QX5I/Psy9uaOBaizuBxPJVhUVA+RRBj0F3qfQ1wieFSB
FBDpjmrwzNdsLhDWEv50tT8rktEoHWx2d5CuV5k+G9UmHDYVlgV4E1iO75M65Z72MKy92Ut3Og0b
dkh7mjNYpoanc0dv3ND9YFepJ2rR5ly+cV8wSnTbJ8aLK3mTBY/O84RczVttD5iVWLPRDFPgCyVH
UY+zke9sXYZgEKFynf5iWxf5GK3hAI9VZzSqMhofv/Eb8SQ1yl3anlTEdaD3BVsc4gowVJX1bJi1
DqtaFxY8UYMWb0Ejs/E9Q3k/ie48CS2hBAho0Nd7ASZnuldAdkEBzvGCehLN9vPkZU478Jy4CWoC
4gppdYI1tzEbANkNJAN8Q6RB7rbEYNXa9JI3lSnbSqaTuDM040cQAjgl42CdqUbNIFhUScizfvMd
kIzi9Upkpv+36VHOsSKY/nsUp9fsSkc4jrYn1RI/zC9CIv3g3OLXvy80DMIoUjqueAAi2rQDPdhZ
82q4BvoxvnYXdYlWO2sPtwYfEuR4BBMFIV0EMqcCUUa0dKGq/Ko/lmo48zXHrVzcWnERPG7BTWCH
X7wa3OiPZ5mK4ycNfQY2j+GpxOGM2HxReH1lPO6xrXhKpIYz/bH1Ip0XEJzXWftwuSh9JpfMbC3Y
0W3MfGcW04NkRUZEHmJojhATt4SirQ0MAEG74wtDC4UkQB/rUDSCs4hG9H50AbiFJyigJoGx7lj+
pVsJs4VszFIQaNUNz5bK1qLv9gGmpZdlaRh7i9MSR1ZCEGzoy67qQHLZ9ApBkOwdNd38ehh3wRKp
YBEEWiPUEznazAmHxYPD+0/XCtYC691aMbXvQ2QzTgl1gZeQa+K3inLowrF+2RBjdJv04MWlrGDt
Rb0SciCHnkv9eGN9jJiwIMuiFS+3yAJ+OaeHnd0AEgeRSnhkGGi+AqK3c0U+90g96RIKTu4J7uVc
TfNtpJyJ9z4hGJQT08J+tQYyepfSbY77NTI915qklz5oyG0WHPyb0aZ7uFZ/yYVeh8bfU7+oMSuh
q8jHz3Dmlu+wx2S275g7Wn2ETZLJGfa5wLvKJdfaluxNHClkClvR4V+EdTL4+tvJnP3uUeGIZZ/M
eb2PKYQT1V8qKKfJuzxNb2dI6lC8HsfDotspA1ppZXse5bP0uqd0FS+0LfyGPSrgZx4kT7r0W2J7
66OREezqV1G7UQ2sNRG19oAnGcwEV3Ny+mgHr+Piv4dDKBB7g0Y16ZWM7uxsfBCIzebAcx29+aXG
j94uI96VUYHF5cTMx6mVStNYMSfYhka7VXC84dKJiGjWH3i7uX/jYVrMB8ZVjboU9kXdq43mnhaO
qx9rKKHhcNYxpAtazAszTf+Edz35cRouJL9OzUif42rhZl+KpKg9rRhbBcdKayWxK3sCtoiuimxO
1A1QfgxYWvAG/a7QfZakj8x7su3VSn2uEE6BrWeTNxUYpxKg1sI4fQFaK6dyneBuE5KJW2OJJqK9
B71kG0X8GDg4+VoH5VMFfEyIaNKgAyL5ASE00X2hWiQ/4xYdDyvhdugvh+qyIdxArl/OP+a9CMZ/
Z75NQ2h78IWWQNmA8G25BKQwYPpvDov9eaZnYkJIMHr3r67gLoNLlZB7MScIVYeY+0+8nrLSBp4l
eE8YwfSgh22Xt2QZsz16GKAejVZccc0eEj5a+LQgEOYj0t6r3s+clhdGrM2hmvDLWG7gETYh82+f
8IAGyFzVUV38Q5aQomlkc/+bDDzx5EPSiVYVSBpc/GGYM4KcF29SWZiltffEhQlNy5eedmvQegjW
H5hOoeCNeuaTcVvRFmHHDSyiLKBrHYRvVftskQulqrXjyHrh5oAp6w/MC8ZBF3qsZ/grieO7bqR+
S5IQs8nR7QGlBM1tzPz0Wk8/eDuw0o4upn/oaQ92o+ZmUD1cZVcEwZEhtqAhR9h6RR7HulSOM5e5
CXVhQZsu+o/vHsCm0xcv3VKDh1FMCmQUSO0+k0G44r1dRuP+uuPukkJhG3FB3CWSQ0iGzLEMuseT
ssYGcGJA/KQTO3AC6gA9xt5aFYqcTHTy/JsyNhP+8QY7EYx16342hYZdP5Ee8S3cGamGOGeriMP/
zOt8mP0txreumswTlZ9c/eewAuFYL5m7iZq1X040l9hDRR7rDjPPadbFg7hskL4K4TP//KcpBYut
oA5uorltXcKXQSMnAqtRyRqYP9ksD4FypPPsIs6ZWtTVL9uxZK/pOK4M2KbpIOSZxEGtR1dokK04
FlywDM1/2hrQDO0kSaPsc2kCGKAbVozm4WS+6OppyyFHt8iDROh5DBUMnerUdOqFfzPLInv+HvYZ
gzOylYRCmFbRuGl4Pe/k4k1zK9L0myxQKHS95vKhV8Ru5mEjL3rJLtcAoWtYm5BW87ui33zjVWEG
iPIzm9+CMcrJb2wayi3GpLoVC762JyfPj7OwJICiLxsioXrwMKK6qtE6lr2lyKRJh0aBIUNzQkQ4
1158b2bs2K1U2kctRGCMjXc+v72AmVLqzYr4LHVkFXoizBL7OSS9GFPWf1VAmZ0x7/IC90vbtfgn
1UNhfmy2zgr3y/a3u3F4m8PFxhRogw63ev8FQoh8L0Z40PPyc2d0ZeBLuOE+jaZVPWH1cKRhWNV9
SlxPWtnAV3zuy764hKwQxYgQJFd7bHw65V5DZ+QgsEiiZZ0Mjda3nGj4oJr9DQGrBw0gcn+FcDgA
PtnxCylBOnJkFoaLJwzlVHCrW0c+VB+oel1SW5byLcdgVrMnpMEdc4DFvt4zqsNxZFbL6EM0wC6y
1g3ZCA2/dP+OFTSadrP3NMMzdkTcOfuPfv4PWZFkcGYOPZCYHRfUkdHSVLRdSh/PDNO4xs3pAfP4
l6gvfAiV70+K+7IMVGAjG28kFWseDLo81b7qCiyc3ANh+IGUiRYW7GCa+bc2bXrNgrf0Y3fOdxop
oX/IndezraG356XFfGEqlMS4R8z+ApBq4byTl/OhjD2RyDaVZVi7B3lr+6OaSU1HFfSiECermFYM
cw0GUS3JTm7QT+7URWk6Zdw0FL9xn3LvpwUa9ZspmVehgmq6ePEeiEvdTCcN3txqSKlRTbOYyQO7
179eoXLUxxKQ9pKk30swDLvJ7BrIQ1Rm3xDyGZ2byiCgG9lyuVeGac37IlQkHobwNiJ0yCY3S78M
y+8vaPx9fYamaRGyj94Fcourus/jly16pFlRO8Tyg/umzi2hgMEcl1Z+R9dW1sw5I6V8/uyQPEUG
rMsl/h8c6hyQYkngXxAC1l2p4/oqDHoz9cTgm7nXtbbL570pCwNd3s104s/xYTzh1PWzxGWEQgPV
pdEBjaDwgy7XhlHqOFR69rtiO9m5VgZ0lmK4x4Nl4wk1YCGZVDi1QdIo2Tj8JU2P74Uz2wVBz5GX
VIrSJakHTidi8pR8vsf/aoSoTT+jEGjnq/G4+UW3Yr1YnLBJFW+IWwyUJONvRIeBFPga6KW19vs5
W6uhVkliIvfayDkEWhP6CqJ38QjtXqwWaWdR1X3hm0aPT4PaVSRca0OidYb0RRlp+RMvFgkQ/VPv
b6ciepJglsItHFmfX0XTSe4r8GxsbD1Jb1BlxemKPyvs0IMOXJl6wfBd0YOpsVXrU6CGsScqrECq
iylZR2SzKJ8O1wE6K3qRd9bkUULSU4wmy6SjVUX0DFVZxlyCy7WtHvYvg7xfM/nKBVdFUjsUIreD
9amuuTl8Dt/1co698udN/4+XzowqKbhUF49MHO0dP314UU+FYbV1TZK0nMBym6m56lMaTuQGT3sG
v/oDlOZutSpFteo5N6mlTF6LFEcBJcqafDgtRymYQSysYw7LBdMoZYz6L5NiWF6M88KjarreR3Ga
9LtPF7hH139tQEzgETdCXNvgDZg8CLDn1brpExZ8LxJqDbOwewiRJMfv7ZqD4qaVxfzDLsn+wI0W
BVVl1///Vo7sso7AZJe1Qg6Hx14ASpEkjdMqQBb0sIEF/WiWu/FndI79hIvAaRPWD6hQ4YqAMwol
9TDIdcy45323IQpt2aUTur4c6XMwPVjsTIXUm9JbdbXKaxFjQaYput5Ti0Lei5qhsO0tVmbfRW4c
NxN/FwQkKMYqfWHW4XiujV5nJcf9LxnFs24oQAXjLQ2IJMbQZRt04+23x/s4ATkN+PDYMxvWuuuk
pCVO+PLMw9awIwFajsrQt9bPSFa7cS40VxAwtc5PHqLjmq9HtuI5f2IL64NpjXCzz+6XoHtn38BT
2drZMsk57fgObGxgPP31MtYTmuAYKxrsuauBsBkwhZTELzBlib2pEyvRhIc1q3F+oq9SUhXyFfrn
f2BVa+NjtRE2eBZF27RqNqiFYXmP4V+VZphCS/FNEee5lLW3nlrer7K+bTxnkRjx2wqZTc0xDmYI
JZY1MF0PGKw++YX2+Cs9JddTtpwxttJevlB1LyTd7AKNEDX5iUfRFvFmOIRuMGMpdqQKzBfcFLNA
gQ/UZP/AM3va4gvrx6Gl8z92aqEBAbb6Vl7eWGwnJjH2etMNvbhTr6OZJ+lmMcK2q67bgA8Kzotb
Cvf8bu/2L87emBOQx7+AQqYUzFIJV2TuxtFj6ic48ZSQTWDqHsmUOn5T8uCemfS8wBFrFAcfDtoY
GtGNleYZ4UXFGQh+u6PqdVhenfijN/5yfxRoYfAs+dVVlSa2T7x+C9YmBPfIv2CgG10H1zCIT7ya
RIWfOB2Saqtfo9J4S3C2ooKwdebf1JNsJT0lAZLBb4vNo0ywUWJHN8BTkS02LP55LCjM2XPI0BEV
XgMneMLh25R9sBgmRCYnXWuY/8d/BTiy/GeqZnhH9Ml0X8iZg22MBP1h/eVf79isufvrSozFodFG
t3iKkyrAr4L94gpvO+sKqlMTbdDqmTFSQPGM6XyJRi01WWkz6sw3GpIxrmzbDsw+GaWFGhV7bgKU
YQoumlr1NY6XqLPzO7U14xuM/jFSQ35RSCljgjl/kzB+aalvNwzHdRh1KcVJUx/6/ZJR+uj3sKfx
u4jSbqUNehJy2z3+byWWVtmlcZQug0G6vkmdcEgt91vX7uL6XB0sl65Kp6FH5lC7MI+XnNMwqahf
0nUMqu248aXd+RfNBIs+tquCQmiBeYzGNJ1GHAiI7iqkE844yhu9PENaIMGmjm/5LYQ9PM6SBBNi
siJ0oLMdYBS9hIF1Z/gsAnAkGre+T/c3OBWEYLUXG4T6FJAOPfs5+lEB8iRbKN58rBplE2fYJTJE
5VrPuMkBiHItTfaZ3OMeW4sAdTknMe0tGB3uqSouWRgGtsJHgZ7E7wgHRZeXlTN/tlgb5sqe4pM6
dIJ7+/5D+0zZMRgdz1XQPqBU/39m0iOZWYbOWn++PBLtKS6kJn/PSlrNygfOScjpDdym/4//KrAW
0vtVHR2upDpj3ZknA5HNxvillIMFYhjf+1wcVM+HYcYKkEU8mFQAAugkCib8/+9s/0NG8bOHjr80
/vQIYy1gh2gfdubiZCCqBd6YBmiZ/jqNvVhryws/1zy5ZNkBkoegtKiIYsXlOAeoTNKuhBYFuBvX
Ce7Jp9Mlp7qhXtAtGUmq2Ow3omQpIfckJPQQHxEHvyvEKFSxiXydrB8yj/jeAH5DceOex8hHdui0
yzCngVp/7PKmODFu0O49QzIXI2uzkNT8k/MarnMrSixYshLX6hY3dku7wm4IKFJR6ziLGp/WYiju
M7mPUKZCwThXgvs5yVg3oYGfz3WemY42vJuXyzU+tIXRCqq55qGzhZ9LGcm3BOVIL7H4FeqYT1o2
1jvNYBbKJet9VmGOnMr41mI15/Dq1/hd9AqCPeq98zsorFxpCKv9/QWJLR2WQ3N2KdHaoBHckavr
W0qNw4HfJxmFrNc9jMEjH9Z2g2A029g0zypqhEzGZWJ3EUepi3KWSKgT3FBaCoAVWeVuyrmFa3QD
aCL9j8HUDIVw81V1qgX6XWWsCnzrfLqpg/A9qlYtmtu6Q3x4HXC3Dyvzx2YQWtB0YgDuYlD9vVaU
zp9I5yHo7TSCOwyeHYSZ8mAqmO4uE+j7AQL100dIFrY3giQH/uJwr4kKEbR6p7hVsFAOgrM9VORs
WKg9I8EpabJ906bfOFJwW0IpCqwezz3bGnqPLUBsn1ZG+vP8Gs4I2+G3JT86l0cV19LRheo8yc6p
j/JGg+ODQVRLvwaSVM10+ZOkCK028tgRlY+J+Vg0x4kF3hyv0O8Nb3KvzOqF5t/GXSw84jw2xP5c
ah42bwFfDwbBDmjyRB6FCorw4e6tbxjHSq0cETkY0alaPq5/Rs3AV4nEbYr+jufkDrLFBLgyrG7l
zUJ3gNVBdUaegLU0/5nB8sSxPNCzC9qub43wYoZW0l71XhrWJi4oYGUrTpEWQv7Qq+b38XJbhpk2
3QtqCpygrP2V0QkbAThMewkZcG3j/mNePmmuAw1VTsmyVXhPdJN8stFQmP2SUn1d++0umBkfm0/M
FtHAZ6MukbqJzpXv5qq3TpUuijvIq/rw3xzWJPEJuVQOrffXMBivUW5WojX9XIS0d1XnIYcw8y3G
cXaCDf2NJMPxMfRX6WOBA+qI2kO/sTDGp7hBntdgdYPEV/mix/h7mX8lgelsCW2BKwr/9bShp777
6mbDfNBdITZG59ghbMpNDR5c0c0aAsqSjkhGYhd74lxkB5u1d7MvZoJMyosf5kSjYtgYBGcN8fMl
tJUKvjyoE+JfwoYuP5JJRZphyIQLrKxLE4XyVWo0OIMuj9m7S398yKw2os0bKYOqzD7gyvGwTmXC
h1mXZaCTmPbA3J90oa0NHSjUx2Pz9gTAo58Mo29wkjlWTxPS6ZD01jVmDFmpSc4tFusAFIRy15ZW
iteNUvSyCYBUu6A8rZtqcMM+YAY7QSnQ5NJd6BLSZw1H6YZ6mwz/QMkaAuq8a9xeLchAOeRYq00c
csrgn++gGpp/v4yKbPQL7eGZe/ZOudJBmGV4Kzt6BETwD8oIwDnPbEAVgUWjx4Pq10/3uS9Dc2Jn
39PnYcyMkPn2N5fnkrLk1iT5dTu5TR0R7SbddOJsX+KHcK0/LG9bx5NG8j98LRp2y69tcqLRByCu
KQi3zkCYQgTbrwT+6Gu3DxBKYKEsKkhyXvzPVDxFAWVDtrc/1wPQq0u7UgxunfIv1Ubn0MbDY+yi
2mjAY9lZXMwRGKka/4U58CWrrLONoka0PiT0N+nudIwTCdFFU8Up2zFCIJ8FFJlgvxLIYUvfQPMD
TFs1meRkNd7ZO56HaTuM4ond4fn3DSnNlK2nf22gsVh8nDeopYP8vC1JS9mRDkJ/rtFhIUnealKn
FWOSaKyMAB3g0Wb/qrksKtwfV18ukMap78mch28y85CZznnBwWwqXEY6EEVxHYxeIz7QYbZjdImv
3FQBxaY9fS/5xz/SJt5jUN3EzHVRqch57MWchbTWk/Of/MWwgEV/CpxGJgJu8XHiZK85e8Tt2ajF
jNN+SBAgabhf6DIY//u2IxwDyzHmY7YgGgjNX2FcrKXa/xqzZ+0aNyOKZ1xlIUOKew/Gwr362cRb
3p9bfALkSFag6EEnYm3UqvduBNs/TWPmiqHxAkyLnDFNyJsoVZlK2+6/AbEpWzgqDDuOd2WfYdBQ
NeQ9ZLjQC5H8SkhkjrGsPQNqMakErqlU3DsJkWNm4gbZ3xMwResAl9iilek59bSzI/xNsjSXMMjO
6WNtXz5xz9b+JWtC2WbGjVdN1cGMWF1tI4Ia6neVgO6yO372w0U5v9n28HBI+WkJkkzm+A8OItuU
CuvxT6nq6N7Fk6WRzJBGbLTYGKuqbmo/oSjkTNkpgb7xN2ZQbezCRbdL5e09PTa7DzXZ8KrtKwg9
EE5CyqKI+5nPEN5n37tsr4l8BEu+J8m+KmPolqfpeoURQsiUX3gOs+YmbQfIlIkzJPB8rdN8u299
JkY/KYvk1XXxFyCgceHPGsq+9IRwVA1uzaq7mTQFSSg0tbHagHwG7fVlOE+9qHTp2RxPyKRPjR9M
DdgQht3INEWf3FquLKBa8UYNHajcclrtUbC2UzooemJIWR2SJIu/yjqQ4wjNpw+UJk6ZDpV7Oeiz
5M4H9LIX2UsjGIWyjy+LMUULZ2IQCfjg2jEiRbMQmAd2ThSBW2fUdr6C/cvdJMcbq7E0IfIzfTRT
tRIl4XHsSTwAAhdJr5oBKXAnN2pKFpIy1LKgX1fiCDkPihSAGi6uHoIJ2WZPCVGlGl7D3zhdhDhH
vU4zlknjuyOZTy09W+FHhWrl2KaRqVZBMvVthHSL/J/Pudg2FrYfY7gWzAgC9ibUMqMCob1Ns7q3
FO+y4dkyQg8xbTv9yp+lkNg2Bkfh7bOw7vSW7iLCy7iD0jQlzjgN4GhQT/E7p4giCC3eWPv0nEyW
57aiibmw0fAD/UJ9Nk1dgkhtTltU0s0EjgiBJFEX+mdb/Qpu/l15tGWCDagGIJaznKpB5+1+jEU0
sooDwevwbneho4NBJTJQncNiAyCBuTtVg827Encyt8Z2LmXldCI/e3fZ7JkL2JbV9zQnHcG8PSQI
0rbc9lYw46cUcopjV7TuIXi1jiSN0lzuMYGTMMPU4orW3FHxj76EpOiRzbGDPh/g2I/rn/+6E7On
5vX7dCbUtWK6lmlWzhHygP1RmypUB/ePLaUUaoLC07HZEmJne2UkNJSqKyICbh5vYsDZuYTlJjSW
sm6pMl3+AcXh7+VYhu3OiXswvz/Ysv4+5fZSVv4b0Z4pJsgrw2UysxLT3aVCywTDSkYBfaKfkpos
CNewU07uWe2rlcffRNU5F1UKO3QeFM7d4/xisUsGh6c4xph8P1geoKHcqwy6sC4bUyDZGeG3LVyN
gIUjWkhUyhS858/AQY+VeyiF/iPjWsvK0qNRYBB7dc6cquj39vhckbBCme1YGOjwYKmloLwInNbi
QYC4fI0JjMb7eIDrChleEZ3TED3eZRhDNzEATeyPiZsPlOIdoKR2eX2wwL1lfcxQNwE51mxOZAtf
e+fJ9brbPSYp00hak7vbXzLWd4dN3AB9fZ0FU6VUq9k/ZzbpGSjKqLATqV/ldnZYDIOob5/fUUh6
OZ7kYvI/eHTdlWl1XgSKiCQ5QqK8CsqcM+aI9sU/XhFwro9PFlvnHeHxgboymRX65w3pf3bAHspW
W23dsBwLVS0LuUmcYTh6+9B6cziM/GO1RXqCHrlnaHn7IyCFsjPX/CZv5jZTEuh+eqfD+ZDM54EF
9oxbbuaWEQUxtpfhrNU+2lBj/fv69cQQstTQN/70d2R9bElw2HJ5B7CkjF7ZrzVazbJQPULm5X6R
FVf2yQQ4zJdJDywEEsQWUyCdA6nd2Bpq/dY2wKD7D9K7bvP5kivSMowbvlWLylPFy0tAEaRkB4dX
qlRBeWVZxYr5zMQfL5ve9yy+cEhhrwrl9C8xB1hRCMu47mjevZpduiQXLQVs8/zxUMDIBzu+//97
2qBze9RGPiktO5ruNNerYu0x7CMWOt4tXQD92CgrvvG9Pj19LeGT6NT5+jJeM1CPsHXXw4uU0PY3
HjcgKmxEsMyMo6NfPJdWSYvwI/zauxScvVZOq05QilKYeWECikhT9Ag8wvuZm+eJpQPyrcxAo4zI
x0ktVxO7sQOVP9cAns77nYwyquxCSLEmWGotyY2JcRX9b2aM4O5+XX/0g0uSvuwIZKvI/z/1ezL7
QFEa2DJo5AqBdwCTqD71sPoucqj9nmSgFvP0USZfludksog6A8TOhyEFXOKDu5viZF3nZ5WTp1fo
HNzMR7vo3rfliCgGmCJQeePzHBYvTMAM79afv6uhYr+SfvZQpEPvhkMXCIw1iiuyIPRbJk1h8MAZ
EoNJMkO+339/pst4+QGBas+AJ9S48+k2igeQ6fSPArALT8qBhUnZKqDIpLvvC3Dwgan7wCda0obs
3WCrMMFNfyyILIRSvoKsUahPG5FtwFh3CYS3e4oEF2Pn+G/V545qAb5r4sx7lFmmE1BYVC7Xsxf4
y2MJCiADFKphrWCYvkt7qlOCwKSsYzde8czi2ppMlWxVNLgtMzUpx8Km4xHQRUuEJwqi2ItOg3Nt
iRlCwKOKB57uSzpD41NKtA22OsMzP2aolti85uwfS5dinIZElVeHDq8CFCyhAdoxdwksY4nyc8rA
8BExVGxn9T0jvb33IVIu8lmQwyAn4i7JbYT0cC5rIwSx5rMH6s7X+wMTrcKLMXTBnGHItOro/Q6y
gk/fNXddXkw3lVTqGzzy+ITixiG2PIDn0zvq7TlQGdfNs6mM8Jda+HtYqYHwSAXATRF5Pl6G+1Of
yxr5E8MPoke8+DN7TnoXoOD825zr+TmJfcPnG26aF0mItnX5GIfr2gCshPEhdXFZrnQknIFaGmBc
sBJGM88Gsl997HvAVdxN3i8IlOnc6ewblKJBZ2u7HG32gPQ3mjVHHNRRWyhIcThjZPbpqxTPOxCk
6XVQSQyoCpbxIKvUE1sUDbaREtTyUeEgPhE7XLHUJfCbzGGbc7wfdDI5A9Sb3jSk6wzZrc2RBZ4i
CwuhnJ7Lc8JiVzQ69Zl+ZyNbmuT6YEXySkIGGrbu7o1xGVUchtVF08VBcsJSYJXG+7eFNvQ67XTV
eLb82qXFarLkMkLJ0rqfcB6zr2kd17LSN7QN2pKQZW7QIFoceJBxBAC/m5eiz5gd2voVvuHk4QiY
8CEa58tLC99G4fTtta1km3VXUMsKw5i1wOMIQ0X5OKkO7DdwkfiVfB7391UZamzzKc2IuGwPgvBx
rdb4r84nD4QKV2a3Jqdf6oJGwTRomNol3of0/1PEzKSKI5WTq+msLsyHFbOv4eww0tXZLFYpQdJQ
wTwwEgND1jY/D9rsJPIfvO38kDSZwt/xviveFHdDzC1qVni3Dgo+ckTlA/CU9jHle+mqrCWjyjf6
SGZjtxdxkBIqYqQirj588HQAknO1btQGElKguJWxP2uSL3AjLkj889VHp8fhr4ibQMt006PhKW8d
nXMSASKIYIkLRsjIV7CGrNCFDyf7LMIxyEyn89lMn/29vJYFwlzWmSZuV4LmQqtZAwXFlWkPcq+Z
HImf2lCZJMdMh2MMCp+8/8n+4zVC1oeSUwD1idsRjssgD+1Dy4qSjpQL4rl8J4oK0CtDrryAbfoG
PGr127C5HxDjctGio1DrjM4V8x5snc+FWnW2nnBgsWAGnE5FTn+7vJ/j/HLywUu9AiYds3wmDPMV
bryLg+XLmePHQom5ZhvXL4U5SUnZ9mH8oWx4qAp5aFpxQlpcJw1PeX0X58ZScM70HrakbE7WKGG4
ZGRXxTMbP/hdxJzZYRwHA4Z6+XQGAhqJUguUsTi+F1yZ4FPhnQYXBzVz7Dl12Fz6ZhCmABcSaF+K
yocwSF9uI+nZpabqD6LFXpEG3lFcEcESdXXvbbBmk5E2Wbsse03dkXo/RopZu7oak3oN4lCAimbw
Rm7eEH7k9+F8NsPsYAq9ylMMPKoS+kQekBor0x4ngwldPZKZutk361JkpQoso2sxgDrqmSWgziaD
Devyan+s0WYgDHyncK3asp3NVM+DvLGKNAvOUgUHAdd2o6FVc4v3h0a0ziShlbGQveKtdSfzIiYx
//M9H9mh4JShJKDrLoBcjB8EaY+rniqcfPDlaWkmJAzzly16ZtRQ4a0qrqFU9EJjyY58aCpdJsmt
Cwncwv7jYh8aEEB/ms5YvNlRL6FTy0DDU4Ud2iOsbVj8DgyITQCtnjEzGFJTj5gQzJ0ConqhCu0y
J/pmFCFpXtwd988Il49tnvQuSL7/VmEBliCR2DnZ7jIoB/IDeaHdLHqSJpt8ApsLw9CfdPYprD9x
FdpgvjwoQl5OWchY+kmVpL7LJz4sReSeUE6lgcF7hqRFEMTT3mQRSbZ+oDM4CV9pMy2aRtLvdfFv
BLI0WjRn6Rsph8f45/lOidJ6TCFH01L6qwaref5L6xjKXxTrN5B4dMupyyBnOlkJaOqNADi8cNCC
Jr8YQGDd+SSkO9pdS0Iqz0A1L+gITjZT6MjXFSkzXZMheLtQLdwlt99owyKTPHbIDdceHsySWtpE
xHGYlh/BuVIz9nsX0rU4iP+19hIeogx/jfOdhjZrpA6xKR8IU0pf1UxYsFqoBDvvi8AmyPeFC8u0
B3BZzZp/4Yi74k9XaOw5tVkValPsH39Oxgk6ngCHZD+1az0ny1W/Hb4+yNe4iHQg7yDvBf42W3wm
8hywXCwm1vBmmZZvz9l9x396OAG02aFW2t27yUzbTaNmeey+MI/tUY/mfb91BENvkJyXJ79rHXrQ
Eu5e0l2ddhfzVorkY/1kAOt46V2ryferWMaCzzE+NAsrNVXqPbChkscgJN3lbmgbuQIB8zUtSjKG
S8oPZfIZaN5egh08sX3pA6QL71eILEGtizfD/64bhYMlXSE7UOU9taKaT+ZDFZW7C/amC3NJBZlQ
34JtaaKYWFcI2ieTsBW2lUQ9ERc8kwKe5eZlm0h4W1u+2Ne3NpkcDa29QAQisBkq9ct2f1SVeiqv
CPWGSQN1q7GJf067BT2B8oSRQG25NMZrsO8YuYJ+r7lj6X4wxtbxYXUecO7pFKejygTH8+QEm9+k
HK+YCllbZYI7P121y2HtePJWa3anQi0FDcGJXpInPQJMBDsPGBqxm1B8r0nNMsr3MzPPYOlBEuiN
FpZSkkrUfPI3FzoiMt11R2lx8zjej5yUfJ9vFy8beNgMyKL+eOX5GyYAcnQ9KNRmIYkv54I31pwR
L5Iaexcqi40t6jNVEXsqjjFI4WKz7kQa6etX39KTKrcn46JhAOHa3gOBz9JaEdQa/BjHnhxIqHsd
GTpUjMS11a3GKj8mvvRs1CxO0rp+PqUPfAVuqskS+x9y6vyMma/Umj0dZqeYmHxbkrMLapuO1+JU
PcG0sEocmXTHnVSn92HisknIEG522cfL+IDAzxKkXWRSAXYuKOT+mPOAEFwzQF+JSdm+hmvK51Qe
R75jg3HVhv0IccovIGjjOJwgOmEuM6TaJZb0KYvTKcRmoew4zrCG66/WdxFyR/lKuuSzzi54Pcs3
tT6AQGu9+83pakOgHXqzKV0wWPRqQL0W1QZwI5+CBT5mFG4gDAzNyrrjUg90klqxvz2Vq5kGl+7R
agvi6DnNyntPzyxWUQx9u+nSOBPJRrssSNSmLYlTfPmKCYBL0KSefCtVqsjdFma6oIe23mlsXfNx
rFxqd+VLWABuZQ019NuSOAXDjMl2hgJSZPJi6i43b8tnAsYDU/2XX9mxdWznkK8ldb/vXcKbqscf
8GK6iyhM4IoglMQQWojiUnRMtthT77K04VKv/vYzm6/5L989YRG6bsOPcUihSSqd9EyDUwP5wVZX
rxB518dmHe2xSzc4uIoriGBjwG7qzPcr9HxJ/itunvvprz3j2YDtHVDIX7YMT6vUJ0t494XSFbbo
Fv8rLrQWezIMwC3n0ZO5AvOrCQw6m2OPs26DxAdyO8cE92vDGZ0zNooOpyvMcf4yMJNciVnMbVqu
r8KCAg7fJkTjy10Ccy0ikYl9p0yBMGth4XaVR+cz9tM7gxC477++GpT50OhUAQKH87AyxM0LBfVr
4fAEST64A8V53a6UUj5m7uJSw4FoSy7JpLJ3FdoiFHb3ZM+VWu9zuMdp4zGAknePHvsDFQZ7fd5A
0hGMF8G22lQdm2+ZW3ipjJJYZfJAIPFA4cFZFC/08+taANx365YM6z1+lX5niQqT2zVv9JXvtWOR
9rC5/ZOgf4eEWrJZFReWf8+FOT0Bim/kd6E2IM61P7O2QSN/13kaOLuEyo4lDAPvqGWOUUDsS9lC
OcC7EIoLJJbNUTctCsk13TQRk3oRQPEadgEcMP7R1gN0jBX5BuFb7F7TUPb22tiNrH2+8dgNkq9Q
mz+BXGPqWiXxGsNGDkw/uSSRNDjBPOSZSn8Nd266ZXZWYQ0dfG84wl5Zh5cG/DGc1x1joYX2e6w3
tczPYNo4ZFcsCNFcoa2g9+iuUjdK5ovNd+26m5vh+JF1CFSy0RdxFOCCRzc+/XgLn5vMu2j0orrF
vIcFXkTlc95X0fbCTo6KLgxvuAgqu8+gu8nX+/vfE0U4ZPKIp3h/xPEIWgdvgYp6177D3ZpgbqTZ
V6znhe3L9EkB8nvtLadzWrbID2T+bkD1tbQWHwTv7BanIPiJAuxtFUvn6RzvHSivPt48kAWMWUxM
tGV01TH5RxQZuKacXXIREY+ABuIxurwBge2kbe3iBCknOWOPwrCLJTQ6h6HmyJnx9WBIaFmFTyic
XjzSlhR5zfWMpRENHXvDRDHZMS5deBgds3Ra2Z80rfHyXM3IYPeEpmtQHMEv3qauaJnjmSyUchw1
ZxWUafKLKQfrnCkxMPbn0K7WvQx97qyYcDBLOdVisVT1D7oRS1ylxmmo1f52CZiX9pOUSvIGq3JX
uxy+4ZE/Un0ZXEDsozc2LYpDzUqc/DUvV2psGXHSZXOf2c7QFJhrUbEBGuadUVYTepW6FwRyn7KE
8AVf/ZlWc9JPP5R1rFBtaCIBKAUiOYWAypgqUA5s6nLprd90IsSWpQkIGCNywlHnycBsxCk5PyrV
OrtY7cAU+oOuaDWgf9QAbsoAP+WfUB2hLBxshtowJkgkiG20HYlmGVaGrwOxdZ0U+BsCyMKWsYcQ
4dKiU33rvnW/c7oF4+Nq4W0U7e5xN4jJhzIeCsWRgpIBWjF1fasojeSIR56ut+yTiQIY+7A4tHx4
6p/Jr+xu8LysBlENk8EOyiaaM43kPVtCHMouLOBZ+x7W4ekZV8YNgykOsuFTKjXSi8iPiK56SgEn
QkmXME1LK9ZuxGv86Fl8605vh9aLdBzDxwzxXwrcsPuyTr2nZbEZTBh/92KzvxQkITF9jAesmAGG
gKwMmUrdsadrR73fC/DdMUiOVCPDIEOCaodfPG/Hq41jimpWAVD/i5YDTYkilRfDxGyF+A/g83R4
tIOmbudp854R6Nn6ixs8TW9NGC3jIQhJQ2KSE36CDS2Bd7/Rx1Yl4EfgaPXJSy0ZeHEMdtGBbrIT
ImVxoMWC9tPVYU4ScD+qpzKHih4I9LEc5zS1Kfl06UDOtdoD7Jxh4sNqHmxejHh2uE3CfQ4rfT/z
xLfXfgi0JoJ5r9sNNPj54Loa+3Hm6oFT6dSNzR2EKIyYgNiupmI/nRshTP37ZBjOomElmi5+E/TE
TonuXuhvDXQ6BPJao2ztAEgCTJ01tQpDwG63FVqmeEm22qFutumStlEk6nYAitGA2EkEeXG+QVmc
h6u1MfTPYpI/px0P55ACPiwDUEya4x+eAvttyJgczhvLHxqlmTBXwsbptCXPc3hfmZASlsGtxHYB
y/ULtj69G+ddc4d4YCSoCjVwci1KFFzbKbuAj92uUw2XcNCHZAYenrK0gBg94RJv3vume2B1C9Hq
z1xvldJhu9N+NP1jPupMppSDoBSyqopWLckqdVvgfD9KzgoOpZjF14Vqar3S0cA94u4pNx73EQn+
yqDs+echcCvbFncd5e+WzjzNhGQHNoHvF82FOY+W/PIes4Lbgj7PnWZLLHarI/jv0EHSikEo4uZK
r2JZPTlKfVZhw+V482gFpJXRnc0vmmTof8KoEafwOc20bpNmiyiSFmX3rhGmW5cyPnfk0L6uTmw3
UDUrA0nQRVkeqLNTAS0UNqgSJAqa8JHjsS3NigNrMWpVLvCRC63e9jkkEPuz5wJQeZyp8Wq7t5cY
9dei5+DZ9APkQXEzWbqWY471nDuknWxd6CbSYsh7wZBwGOYfkpmHvWLkC0osmSNVELLElfs8xCFi
MKwpsjCyw3Bdm+ATCx19bNPie7Kqz1O5BEh2jCN26Rb67TtzaWN4m0VV02HixrDNtG0zdN60l69j
VDlZwoh0v+O4om2BKOWsOtI4rKSl59qLPMTEU/S+2tv4E3ob8//UovHPu6TsEm2/wwv76OuIEFc/
NqHvIvQbyRm8U9KJP06cDoXNB1AUF2Xx2WJ22I/RVbVAC+c1jyTWZVGVgL8fAN6QIsE2I3wHR+cB
JX7R0JCfmX68FEc2OA7fYPt+Fl1/yIjWEQ/fYeqG1QbdZyRwpAQfseZYgQdgPwb62mS6ZyXoK0tu
JM9g5RJDZ8eRxU28x80v29ZbPhvpoB/OV7aG1X5hoYIOUCj/QhcPCNHGNP3P/HHZC0nmQishphHS
GOdwE+qLk555BKanKk6c2aBdcZlVXOksjXzIN0ioDxtumvNiG2VfhGZqjbmINqtpJPM+vgPgv+R4
5Fr46WABc/ENftWIjKbi2Nxf7/u4PD35K0xKvHIlaaY4Z90cBrALEk9OYp5QjFGGkxMlTZRZKTdd
zaRktBSpE4iZAF1MRZsvVfDOsQ6q1ebAWpVDpYln++TCf4DOF0KTXqRpzVfq6PE+nXRMwz1CuFtu
qhB/fV6xyrcZEpHMGgXTtDLyPnGwDa5M/jeWO2ZtZNVe4o0Znb2aXo+SfrqG0xEOus2Q/SaURBA0
HtVCtJmFuOxHcoL/La2QIEgISmK1JPa4Qv8/6v87YTuy4Sq2fTjULPLUIkowDx4FaMOi5ldQGhE0
hQoE67356HnkDj18vOeE3McpPGoOVVHoS640wL3ycml28AiqYB4LUrPxseSu63nRk+pDwzSy/jGk
bKdsz2f2jlHtb5rM/w7c69vEppBvZc5XiNad6y6hy48mlfFYVSynLF3dEBK8t9nNDVzmSAyOOjqO
i2EIDwPrqEadTdR1zDKmf5Ut+rdDJJPV3GFkhH303sw2pLxGeDT0OJhPCzExdyzyyuSZCNkxMG9R
i8LxkxUHqFJvwwBRNp3cKDmdMHb6/PhVthlXrOQAsD5nAFlKSa4GE6Lxwf/rd7KnchyvxuOQdzfA
o3Kv7MSOhHgA5gFflrM6NMzZnd09/RQbboulMaBlkt9xXDkld+MCCUK/VQREh9NdJhzDU0BwwRH7
97ozfKqIA/PswwtBoyfETkCJOh/Kuz3sAn+rQGLfd80QcoPstxVDwOlJghabhnrLFywTsVcUL2A1
gjtvy+WF7a7nNI1oOgNgKQOBbDU2MUbjDyCivlw4A3RrVaPhG8nQqKwdCEBmODwnbmO9FgfgTWXP
MYgdL2+3JmaqKISx90XpvB1c+SvYKsh1CXx4crWN58xG8cetUdyaBL0eSsDBz6KF4pfeImc6cx6R
kwpZo723WOS2iAEojuQw3VLRhVv6ji8tbpMgURE/91JenVmQvaPRaRsg6V/mmr5KMEXKQqutWfWV
I+H0IWoB5dVdSNIReakQPvjyCwQ1DnY/UoW4HPYp2mrd4btp7gpW3e6p+JxLJbIpLwajvXSn16gR
n3ew5WP7mCazx/Iq5MQlCaM7XLeJmcqlYpy2kgyXp+NsXyDmuRlDhWwE94cATH5MX94VXSgIuggT
bZPLuEss1GHXWx88hbqDuEvRo4SKx1BcBFd10pln1aoJMBqCYMe6fvCSFV/bakzifqHRiqMLGvU5
KV7pDJDyXx2hntIVJ84MTTnSSlKRTa7JDOZow5aYtCKo7AbsxVct8f1LZejbL+0BfYqWIBf2bypF
/WBGovoSAm6wYES0yRHl7YNwl5QMiOYHDIOtNKtR5jkDRn6HUxRl0GXiHaq/K/jyC15h4eQKQKBk
D3n1pGUgtdjx3pL8PViM89Tzr16QyYeoqDqSlG5aCOBlJ3O+3xFONfsFlcLZ5jN4qpjTOsKKotjO
bGRWWx2CRDjv9iOVf+YbSPI0AA7y9ii+NfAzIke6wXnIIfrfwg/1MXnUOV0de/Bk3cjYSuUc4Jed
LYG/kwhwe9sKod9UDrLDc9M4JdE8a2Y/ThqN4bv29w/JMXgdiebaXCHVBrVEpwK9W41h+mP3oWcA
mgKcV39soaCL3o/iYn6P1CeQ0fKNM1I2wxvEEhGKrfSFBg2LJU6nqXt5sl/SolRYDmBxfxE6UO+M
Iyd0FINKdnY+KRL4MhcWrqsgVmdLCIs4gGc9/YZLjtaZB5D4oILrFxwOMZiFzqPAP82BfpQWTI9d
juFjOPuVTrr9iVGwL5/VqHNFRhsRXpk+NBS/96vlSF6NLyNw1NAmCr5DpzP7vEiTB+Xqil1ZtNeE
1EH41EemV94K9GeLjfqZFVWxyaDVPBl34jSRs87/08YVehy9kz0wSeQQDHYM4BqyYXTKXUwJz3Z+
BB8BKwU9HlH4XlRQyTwGiTw5aKNSNUhxNQlVzdappPyS35IlUUTo10KdajvYWjJQaZK2+tvyUpCj
ywjAA5Sl8KRj8itu4Sdl6I4iqi0ql1VDHi5nVnynYY94kd3HXdX9WmIKyOJ8W1NYVG4oHigLOEK+
Rxdh8soIazSk/ohdlNnCHs/OUa0uzY8ZBrxpi2tpGVlmzfXjkVIM262qHC0BLw/Qq5Wbc1KtgwOJ
tkmBPYmFGYiMZPoNIaYjjMWm4y8TI9NsmbiGCFpVc9U/OEoE3IRky3kfbnn3bY/tc92pYTF/Zp63
dRLcqnm8q1NYAYPej0F5eKBeFrahwfz+d1GaRyhjpB9GD+mBB31VdA3kVIxoy73R0rWCmBHmGUmu
BkttWnbT+WxbHNrj7NbiFd8irTt/UqE9/bwEwLaFHFV8BqA+8i6JdNiymMFe/iwVZtD2kBnC4I1M
FWubtib7CVq56g0CKihyIWg33E9g5vXPyUtRiSO8Mag50zzwbWCWZKJGgiMddi5ek500QotTipZl
z9TtIVtcV37yUJXlHLFFDqY0CliGeVCYlGWWSfND8A3fDQhjnxlHHmbPglL6zURmVRtj9CrHtyWO
BzJBvw72pBxILuE/ZNXn3W8b7lzOUrVyaUHzgsuR0Fe9Ec8EkqsQcI5lFTWsLkVn2HipZsppUwMY
54rDJQGy45CIA0tnjBjwPh/jtV7K1VVqN42CmUX1K7p4x+y0YhWSQtPEn8Q7+/O8LZ0ITciVIntR
HWgLiYLZAgEwBprwOM4wZW26NwRC1OcR89+gAJbD8iqmgXDVqWxv9WC+7I0NxT230hJndaJYgu/D
+RSJC/t3qdsGEZjLyOsho4ThpaOHuTmQIeJ+XH75+Wnnd9CSlJJE/E57r3B8dkF/L7foJMB1+KtJ
rxzs8/Kx4WXLD0fKntSFR2dXQoO/N5cHteDigKOtA3BLlXUNmD7OJDvCmXkYv0uiP9wMOjNm4Z0F
NJSSb753g7ye8TlLuamUJcfBWEUA2lrcKipBjEVrGrbhfFNSoo60ntE1AgllzAfu9oWy62RjOp63
KmKWEUqkE/F0Wg0xs1Rfwh4wHlQT3e1UoQft0yp38nhlYGXUY1pwe0ZBdlUWEYqcDAMByltmwkZo
jR7cwxVIMuBeNg1fazM9uPSmm8TAy1P9zrq7qVKkgBcxPWNzrXsvih9Eeso9h020ObptEGRz+l1F
Z1MqLBpVPpcEvcoiOn0LW3u5kY1qoURvfvI8jwc9a0f7jKDj9Nvo0Lo1SKb7FFGS2a5WKEdANGhM
GtslL+wVOAPpxC1ohxXOCczzU1QZqbAmvDEMp170XlqW2ZTkqEY8Uc4TYiDtju/Covaq/VMUniFz
UIUcrrAljQEwWll9FZ0WilZeLxr12Tw+GtJxSscrlFb5Oe6NOKR/K7e20baa2DKE9L2HAHKKrDCn
IFFheHTVkPKi4ImV7YE7qmp25Ln69uqoHj+DdG4s4bsT9S158tcaC+wnppLntmcafOZU1w1hlD2q
+xvZqzEmyVbOXCTd79fUzkbGGz5plTXZSTC1yo9VNX56bjzUF0X/t/0aBPbK8AU9i5mRuY+TGI0h
VpxjnPGloMH8LV8mOrpW3YTlisXWAxBWezbCXo7KqJb0jDXfzXtePxW+1f+JYJoJVrIkvX7JaRcH
3xe80bdcklU0m7UUtvY5GTPsRcmzJbplNhUPVvGPZA3KDPUhKSTUHjBgPaWwENF85kDaaCgRslyr
E6iSepG7Ec2SA8kp8KE6qQixZnO+bBkYbkWT08gukYX2FqZghZd51x19RsUcKKnukW7E5YQpBpz/
YHU7fF+pHZkUt4SWhw8FvqdcKDFwjk4VEVBKn2iYToeEWQx18WoaBjyVm002S1Z5LjoccEm5ke54
Bcp3EXQl6NMIC8rapwR+jfJZwfni2a1QOLnwqYdViffXdYOGnZ9sIDXQDDhPEmLdAbNQRzCEj6aM
AyIsLwvJ2aUt/1nkn1jXwjDF5xVBZnF3HKOx5Oh21bEI9oaKzOzkC/RI3755JL7oSWz4E+YIw36Y
ljJDl/5y+4C+PTBhMJO7K5gvob0ytvUJhdoCUHZk6N3x8wl8ZJfpv1bRbTLwPb0jG9nMieY2dNBf
/OiG4VZgLjjuvu4JvZjDBmc9nlpjeeTyUEWUVGy+ua6n18SfoFrM7ISq9xgUzTwETFoOlrRqEngg
HzL7ZfXuLALNwVBuOmFrs24qU9qNKFiBddlU4uelo8KuJSJtrOXSLxNfOuqPQYzLzQY+Dxfg1lZQ
+82r11a7FBojomJ1Km4b2MIae4ToOGkXwuSKjBmXKoYAV+MxQc3JXdO2ZSB+wipG/8iduRF92/A6
msde68+zoQScqKT/R3Zsw18RkbZvmk8oRn2WbHtbAPJVG2P443mIikAY4FY/Xj/tE2I+2TzE6M6S
vaZfO5W7f2Z6L+JxpLNcWTcB2XSuAYne/DuINzAlq7guijbVJgMfDc40WzXdj2EjR58RCBt4B4PT
JaKpPh69vrLiF4wCKl/LsVhjldTIbQMD0kuFUnhYel5iw9S0Slo3C471FHH8It2WsqrEpe+jqnym
hHmgjf/ss7/vC8X83b2ew/oH
`protect end_protected
