`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
gtr2VyIfBPHscysZZ6sBs9u2ceVcJP/BwXEisWJerQu7ngAL8H9uO0B3b/e4vn4F//i02JqWXJfU
n9y7sU5cVQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pOKYRUUuretbS1ZgPk4jfRtKqbEjMeSl6Zst/lGM6ZdE6ROa6Zs+W980T+i2R+HjD80boJ3A8J08
QdcVc6U29jxpbzMOz122JeFu9q83to2PxPPBmzaJQdqtiFssddD/LAH2v7kBHxRP6fzwDHL+3ivO
jYd+ZuTEJNddh5XcJtI=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BHLI4h2+GmYdBQa2swfm9UYT7JRECiq2BSQiAVUMYfLnDuTMtIKSbfxoOK/n+k/Jr2JyQ328JGBD
bcs87MQZD+nSVBF04g871L7D2sVB/voex5OvwOSSIHHROkVuASqDIYZh5aXIu/rvFHujQCPO+Hb1
btnLh1/WjAZPx+x3TkudvjF6kDfb+YGgD8gj0IcjGWftncYEkSJWgoW53CUGX+qks/pdzESAIb1X
2qsptxN6nP750uwWKE/1Rr35+W+RDB6MCco2d6RXznDQz2U1Z5mKjz+ir70+bENFg0XH35feMx4s
l59YREQCe6KzAwn1+0gRW4cYwm6TfF3sUMnnow==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aaQbWweXBGW+gZPXQn7VrnpUQm3Zke8xnMxKsYMFqTb9skSrTdc5BAiAw5ygfQfzkxMBJZ2hzCQv
w00WcyjQQ4nZd5x6Nc8bV8q0AHphUspuPatDsgvUYC56SVQd5sZYRDFi1rki6ZFmgxcaUgpulJit
By+fPWJuWiT+ixWxlA4=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TIQhHwMNfE2Na7ADVRCsVjpaslLxz/5GARHTNCio1sH0MrnqSrtDwMmrhFHaW/8xc43AqpwqoFvR
xPXEMmU0y/ykLPWpkp4fEtvnWyibd4VawgPlyjbVsQfSHsfW1UeEqj0737kKqsWgY1DzbUH6dnhK
ry/8oK73v2YHKuVAwqxN97uJ6Si+SmJfqz49/wscqPCVWLjZvoGPZ2AzcQrcmTGyr9e/1z7ik6/p
nm/b4F26WLoWga64te2t+gVIyuwsqtyov/sl5qF37jjwmyoeozbS6IjXXeZEeMhAZelmyAtKkNKP
Ft4iojFLz3P7g7p6WgXi1KL57UoauzIwIFkhrw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39152)
`protect data_block
VVmYeOOG266A8tSL6Q/Izuv9IogMiiUqBsziqV5BpLEKMkp/xYnwXdsJgEnEW8dkFHbClIYukN82
Ds8eXmgwlQ7pkQW7vsv1rs4ZQ5G1Dws6eNeIVEy8ygp+YUz+tD0nY+O6o1VqZ+qfzs1/5Wz+F4R7
HjGPzVbSbNtVFbBsOH7U7Nt/yVT314nVG7u5j3Ll/Wo5AGEyNaaRaQdoxBkr/I34v9/vRgxxHCf9
k7cNqKl+E+zDyFjvI2HzRYMz24PpIc2rbcXNNzYWDFyrBBEj73leETkb2FoV8jHoDEhYiBZDiTv3
umAHZ5kqmcsHrs0XYgVjrt/20hzbvLNSIro8vT6a56F5E2sRHToAXchhQ/MkNsyCLGDOv/eon2r/
ZklKsuG/4LCumwyxak5qZkDELIk5Ej+vatO+YhYMBXYHENnj+CU90eflOB6gYcAJx1+TPbdGFmCD
x4nkyeVGhQ86UiLsXcM6bVMcBkS01IH81MpkscW2+XwTdm8DGFBXBeUXmKcETbWagi4fZQU+53r7
3JGcYa+DT+oTQJaOQzWDIRLNfM9P7tNcS58dNv5IKc9XJ/lr1ckWDT9zBFKHxeeKZ15vIAM2Thfz
52pp7VJBg4a075a/ZguZ6PhQepn1ykh/hPUuzNEF+/8Pcs57GvixvL7XWReaOnn0ofUeNGoKp7gV
BdSLAltDsiEA7vA+Hi2HayB7pAuVlm1yy+a5xzaMhqIuujPo/EtnMQLZpGndVnVOW8WQcTdeD746
dp861LPHdsdjKrzsgZdU0PwmcCukbhmmrKxr/hZ1fNbNIL4Bktasn5PSxZtuFwvqo08ORLcY9z0H
faWp6qNdGf2ZLZRZTDRoQs4FbEb0gSC49PLlW7TFNR+L6GAljmigKs1N9/q8U5GCaIXNMKIUgyai
7jPS477OuP4rnG/KbupxEM5lQglZjYKv4Dy9cDX+B8TtPVHApKhVoIZzKXnf7W66ItcKtfeMrsrr
DnpdFF5VNv4iwuO0HKiJ1yOQt+8oHnl2I/YGcXfMyJk0YPueH5XFVEr3YUI2wdtG+U3icWQnIV/W
kK7y1UJcHf74RoiwX7/M34P1EKe+66AqFluPROkToTE7vVeywYN4wT7XKkXsuxXBDqszF/O27KNr
VzWEr0ypNYDlMwAm4WM2QYDNXuMnl8ExgXvbTOh0FAnKHZNuG4n0p8FccsfppYIP+2oOWj8OeUli
JV/xsLj/CyjsMsHOLq5kOjCrf7vjRqDmOMuRoLp/iDrYWwUqcQXAeF9HNvTUCVua9XA4NmMiBAci
iFjqtsH2NrDnY44rUo3CoUzX6hb4yI3TViZSBEp2oei6NrbygoCXhJI0UFNvLyl49kO5OXZJ5NaO
pPg/nY2ghyEZtig0luF8u/+gvA2dJK1dGna63MVBH/bs6Xfk4DXVG64VLWMaiwJH1szhL8FGMldv
aa7nWh8nfzCI1J9/0kGKP4G5orYX0h6LsYaE9j0Q8tVuTr73aXdUBoSO2YRCP3k433RjYTn2gIXx
FiAkowMnFkPq7f2y7l6uVlHYb6qulXTnaeonXVf8q8BiedxR46psUKjeDGG0neM2Ay8uq2D+1bOY
mbprgMvmcLLMWMJEe9ppRra+SxLGAghSH3CKGK3DQsR99AhUUqWWmRcK3aPhJZmb34qULz6rj71+
f11SZSoSRVP1XlokhLSM+9cTRGKM7hvjrHN1Ps8Uy28fEj3rnKZuLVabsH2gdDbzRWUgP7WxmiwK
8Lds14RFzMatjKcz4IYV73mJSPFboXF68Vmr6PWydcLN4vS5FnEzsRnl3PLD28M/IeKRJ8upTwYX
6yXFEJA4dTuIrno9iPvf6TtKoJVjFnbQaE9WRGulE5uR9/+imqgn2e23ZLYZeYkL5JTnZDYhgcUn
tiiw6B3UcKLRaIoPQagAmPK8zUArnM5TkIg5pYJJO5jTzwRPRAw/Nw+FPSFhcbgevlHDS+GFKn6o
oN8Kyprwlc+J9lfV8OzsaG4e0Z6d+fCyOI/rGIYjiUGcrqKSrfgl57jB0C60bDYmPwYX8/CDW9tv
exs2/gj1GquGNUWQdZTh7iNo2QaTODcSryTgA5YE9Pg7Au1OJSCk+EHivU+Mx7GIQgljcs22JPEx
ame7TWVXgrtD8wlFarmaX/FN2Y1IuFdn1QYxPXbaxKG/HXabKEoV35eme3MqOLKKWtSoH5guwDDY
UwNgklCCidZljcSXCJUnmQoDgzzIu+OvI6gLrrvuvgZQkpxCkQpzOJavGcMLdgU4NB7NhEj3YiLM
AwR5b1SW0YRVfLg2ZzyJ7lMl/lNO3C8Y0rcDeytmlVDdDEc0F8XEUAnV8DQuzLYJwU+OOBfJaKXk
aIuUMpTXrq4GoJpDylFvX/r1iFpjtQMtlvWICqD2zqKk5GzZ/h+Cr1YN/sOVrbnFPZhI3owlsZhr
P3RJQjkrzw5/+2obH6N7a3sSMnsVzwPNUHuA13SGmpL4v6blZHrxPxNFa0EjpU2sfcFerK5pDAkt
f9/XjAbwSvCZKxesUyJjN6bUXYTzxAsYQi/rxR9RxM61qgLr7uSq8LdgHkqoDiPJTmrP6C+rqDsB
RGnhwajIEcV0xkVpW00BzApQdKOIZiXcL8upzmVJPOBhmiMkid6FEuhdXdx7ZnxhYmE36RXQ/OG7
RFUrI3Dc+gIdzAs38vKOmXKn9XyuRWoPPltqXrD6pcRA8c88oYSO1oLvILr57cEbwjqWYVmsPuRx
vlRP4D7xjlqn2abl4m3kDpQQSFB7L1G8q1/GASG0as19aK2i1Lq9lsOtMungW9azkiOwhFO0hVRS
FOehigoLMdCmGollb2qvZQiCFIbP9OYys8j096cOsV3wo5VMszVE9EIsbgEQ4mzitTJkmpJjABUI
Xq2DrDcDgElGZ8QxmJqfqQt4NutjFHSiyeB8VkrEY231hhcrhUSxDB36JZ8dSX0V2MGpBhqemSRc
rZREfSQRfBp7biVPcX2NnsqB8nt8vhmGSlTFYD3Po5y1HeHj9kboPvlq8hWuNcAnEEp+fEWMcFl5
tuXJCkNAKAeovqOmIVqdv0jVzG7qLgfKK7bBLTL3zMm49QnqxDEzuN0HwfNvsjCeQVzW3pqn0GlX
0mIWrYx3ZPUYjzcyw61ZW1lh7+9GVnPd1VG8BMtdHteIwUJkiG14cC8UVNp6ZOSGnD9dODE5Av7Y
aZWHrAANHUAlQ2D3Oh6+3tWiYmiUpxBBwigKVfQ8ubyV+yFdEc0tDqwt10c9TSE5BvzdjH5PKGBp
p9l1SqESB9mny8NNBYCoa5Z6f4SAuO2BlC183Xc1Z+dgj2mb6v/Qtel1kxcJeuuYbE7PjX4dzyjp
Lro5C/ucUz3g41ycBnXXobeLonbTOPnENj/XmZZZPst8YoTs6/78Hz6dFYcpQLNmWftZ5i7ngW95
+2pM2XDAs7HYsTDWja1g6clyAxTADMW1vZlFr1U7+mQ0sSzEUO/3NMyF3Y1w5FSFFO1A8gsQBFul
MgfcFmr3l6PMyY7nLDcZObNksH/R7UJgRf+7hquhKC47gYx5PdP04TQggkuRA6bGk/sBeGSRLiIm
SbpYi+uo69J+AXXI3CFQ8Dql/0AFrAogIWzS2QbowuiZNcinYfXUme15kLHYDq2R+gjkX9AYHgiS
HVsr6HFQQlqTsNBxnMHhroNE0LYpc8RYwdLT2thpoiUxkTGCDQLYSSr4bEcM8xiUU1uBhiUW7Gi8
dAb+ImRHwOK+0v4MouoYFhdTU7opVQZlw/bSW2YQzAtW/WW2gxpuqbYZDK3tI4p1v162ubLhoSx+
+K2RJ9CJZcpvsy+HpSLVFuafkLLFraCtu3VDJI3uZtkhu1RJteYA3aTY7YjTv2UWL6sgeIcmzvk7
cYM8pady6vSCsN0OzpgB1Xn64v3F/EguPxCF8JBHHesUxcMQe2ZUq5vlDsN0Ub3yYRXAuEieKQ1+
ypFCFDONUG6T/CSfkau+3yiUwxDGGDLNoErgC/8FDhR1trWLx0ToYYWN3SzTDZJAV0XiUgCdNocy
TClxk/tibfHYlv++xVttXo75h1XweN4v/ZraS2RvD7kmsS6hCiqckwPCMCo76yvqDlx/RHG41M+Z
Z1rqmMDc2oxtbpW/KQdJGVpyqqTR1O8ae0XQPBHPezF75Gh73afv9WcesMTBOSpb7B327I4E0ebD
VLXELNOtkLLdN/9YxnDg13SVuMrEOk5AhQ+NUZoYg4lsEMYqSPfpOnkdTZZ9Z2VRegUNVahWaThH
YiqAhkd3NUDgyauK2Ca1vUEdf5FcUeP0zcR7w+nf22nvIzXPIKC0weM6RiwP30oUS1+K0uCi0P6p
ows6QM07bOv2EKVobUSI9/ODfO7j+Bc+nz72YQnKVDgc2kxJY+40owyc3RQwQSkEjMDPGCKQng/S
mzvkeJnx8Rz75Z2Ak3Gi8muma2oeDePBjcOvLSI6MSaN2Xrg89FCgpZwwbB23EA4eGeGgQX7sW92
6wcfUSgvOHDddHvqL2pzjvomoZmezuyoUQ0sShcMY2bREaeS872ayB1UxUmh3ugu/MTbC6uwI7lE
SV0fG9jRMK/B6RfdZ3xVSRteFh3cc9sU52KzufGm0N5Jj3a+rKpRU8Nv77LtRdymTXdxfsw13Ssf
irsxx27nplX3TVr8JkKPI+CUTqiU5fBLc2bgk63c1voBhsT/toDEyRovdpzceMXBYs2eCS6wg7ys
j8n6jsA5kQXGxSmN3bWR1obhUCNP+mz93tzoCQ4i+oN8khcvsGi6VTbpP7+k1yTdPvnPVBESyrI9
jwT2dFv+KeOFR33qpNlzRC4HixqTHG2sLznsxitcagrnMJWaCjqqDfBW4VxWta4WA3bIOQxNiKCT
iy+dQT7//+arzcfnonwPDgERuUGwfKoyIa3U6616jwvHJV3KJSZstNwu/zkPRK9ZYIXGKMq6gQkz
HY3iazDp5W4gMStagfceaN2HxYAjU4PWSTkoo4o1C4NUDdx1VeJqQ0iiKsPDIzNup5LSefYEWZBd
zqV04LSF4MkyGC/bU2KRxYpgEszyNz3RfgW2jlfpJqqq2mParW6voUQgjjtKWnQXmT6esrIpwNVT
uOofeh8VxmTIlCFfFPDRdCf4q4Qn0pmDnsKjk+eKYU25TLcnG9r69VYKtobTbsTUBNW0+PzYHGZH
qsaAULyet3MTeV1qHIkcynvU7JmevsCyRQPhDpTnn9U3zxlom74WtnnusDWYlrMXbpaEfG32qlJN
fcJWyUzAxm2K7uKgGmZaNWm5v1TE8GM32aqhI0JZYqKoTMx7HxiynQqTqwQJ3H31wlcCGZmJxVXE
BUHiYin4jz8hPhBGdhOKU9VJkb9gpxuEz4r8bjBHuNuUj5uiXl+Xm7avqTIADogQ/MsYmhBmBL6G
TnejD5KLR7w/TYLsDNRPi8zIiFJed6/UHfv5cZvJaFXJvXJETY15nxbxDs+5hNhLuayv3gtGu0zZ
rnXw5lkPd/CczApEY76CZyvFVJDMu1KL0PFRShl5si7NYDYbU/ImkqBjJ6DmLxN8sm0Uw5W5uSkC
QQ3nL4LftIZZhnxhlRpjvg2jFEyu559c29zke1NxcdSxLIoZECoVrCQh+rsy5nnh7XpAujezMkUC
vSHSXDzG6eXmjI4BUm1w1o037rdVEHHqNe1wKhkgW8HjdleEk7KjkJVpKTTE3m3fA5TrqcdUv44h
HPXojtTgCSzHa6YRH/4aPdeAuD3DM1abvc6zjVLQ7lfHhPbe93q8VYAw3qpSJ8YBByWpobYy2G/7
eL+O98V3IBXm0L+7FQqGt8GEnvLOhQHnVgNpuVea1hRgZnxB1uSzKrimRcz6MgiGMbNADAlDKP2e
ysQ00QMrepvAsMwxzb4VXuDuCzv1BWZ0ZrICRpwTAC0iYvUvzjlU5DILm9GSBro4Ln13/VgqGquM
Kq/YU0cjfPC4+vpUsgJK2BSbCgM1oPvQWqJfoMsUuECEIr4brQbSx+LKhUT9KYgr5qo1FJTXz4mI
2WUYl8ez2rbgSNZguf82qZESO7OqxPI3Hi4cZLqoSj6CQS8tQsjnozwSnQh4vUfh3K0fVdP4hzVW
rqHT/8EA6cZ6cU6fYg2g9m0V3q0HcC7IxcvU3/BcHVDlQ3tAnNofoaKbYuM39fyILYiJDHMZEV/d
Pmd9yqJ56MA9ez0aUSBw6/c4EGO8pPOV1BWxe+lJp5xUYudDcm3bw8QhZRaqoLfE+/dI/s+TNN6P
1gYKbgKuxem8AnoiBRBnKHKzBa+gG64oPVo7GNCyfiB6j7XqJRvmHKnNu+SKDbK2Qsis3cAXWj32
4NfRaAGu4hWnekXemYCEJ+mR+HOoZmvc4jW+24AU++8KDMLq+cKVef6c+1AyqnSbnXl/ESomM1hS
xJgyx4PsLe8u/8xMNdy9HTADxuojtmsZFepBob5Ji+EXGHrEnhFwfMzLredwVqoy5TQCN//+AzYb
9o0fq2q2ycTCncHoIFBbgElRa/2/pD98w9Z/sJUvHG3orQO/akDYLo4UHEY+7mc/4M6FuUyKyciu
xC+liTd5Xcg59zu+R7Sqx/6utqU1QxQ2KYqx9YuT9XcgPCCE7KZEqAm1gGkwIcuY+Ux9hw8MXXMP
TSgAddgVGJzM2tE/y3RQvxQ33yuqPwCeM/JKn62Sdq01ItUMWVLdlvyCIGbiVt9OIijkjfE/PvNj
4Ss+vIdcUkzAhAUSe/7sYLfQ5F99unoh3fpJWJID92n/Fqne0lxdycBBd2sJtG+8YlmcWKbUkhj+
vlLDZYSPN7AndxKrIqzd6wU24Uszw3rN6gc4oEYAEenRcj8r1qIIeKZW9xo7yXsxbhKMcxRFuagH
QG86y0pIltwby1bXWWWv2u/VaYvUtkxlTMMyFknFBY4ehIhZM1TAiFWegUJcTsWswjVT3h4WRktx
vgYWTWWxzKUut37IsvImAyMMlN/TDADBzrsX2EiI4GbbreCwp3MlgvEys4QgBAVDRbehQS/euVHB
0Us5RZ54zkTBvwx3EAj62PJcEYjPFwBDYy9ZxsBvT3O2vF103A7A6OZoUzIqDKGihg1/Kz6Ur9y2
ZOBDWfZFu7DpqtDw8GlRIvFoXdXUsTvwDc8U94bAk1mBxapjokmEJVrLafWWwhE+jCrskl8+UHzE
pvQbrodeVLPfe/vU39yn1133lDRTYw8pJjaDkz2OoxK3rOaEL45G/2tHoWtyJMORx2qnMRZN+rAp
V23MPvp1RljtFuWNAGU24gN+owEskLkARBOhiJZIpj6aq6O/feWwpQhFiJxcLjSD9vzc1tvDg7Pr
2NabqwaOt1mTu2WxK8lI1qPlAorvv4GioM9EpiRbQPyx4nBAhMGom8OM54QUPzOUNHfw/8Y8vMGX
c5UvnBFl36Le4l5RZb4bYIzuuCKWmrH/voaazfRQEto5biZ3iuwOxY29xc5vb4Ap0FIMyruvmNfI
AzpU3Cw/CDOdcHqd6fnXfJizAdxpO6bOFYHxfMt7xsAkUCNs+v5JoA8Wgfi5rp3wmB6odFlqUkka
w6u90w+/Q13lNHwuovhgq7rNHAdzzJ3eyzL8dEKK9U/DrPhj5XOJgNTGFjlMLJSKKhTkN+ZPK7yK
G/BZ/NKocFCFOAbbPJ4wQO/LamEAmnk/hyURjsfNWGE5vlxkw+wNg3rBKIu329SOVfu8DITNzEse
12eH7bDxLaD0+fK9jOThJbSolZJkRK4T8ELmkFswHcIlKbXbi2jyO6OkOZFaDbH2jJdfgO5H0mb9
WWdCUChuMcpTot6eR5oUpO5rBWDSVXCAWLiKvaxlqmMceR28mxK8W0KzyY+69+AjngRy1wd8Bour
Skxmus3vR3R4N2CeboorbqQ1jCnafi/y52Ed/vo6ttP3eFiiuINb9mEJofSHNM8HtD3jBi4jGr39
so2gVCTuWzyrHlGJS+2erl2AYiN6rgAhHUTnrXGY7a79EMCz/bbaF+cIn7lOnZXC0OLXcUL65Duf
BmvyWtf4n26YI9fPtjuTUmGucHw6R7X+1iaaPGSne7h9OcrBeSdlKe9och6jEHTlKqfaMI2OP1ug
iqGGMdyI/w5IcXlJ0QoecUf2/mcRgUSB5HxTx6w4bD47nMAMGxysCcE+HtN0I4oh2kfzHFwvg/vk
S7DPMf/R5htAA5VAVxusA3D9PaZfi8uUSSisYBahZdHhVc9qQljtYxDQbaqGJanDMeQKQzFC6dFJ
2cNFk5wJBp/wFWIXyN2+JbjMSvfqNiQyyFLA9EdMBtv8HOTZRRGmlTQ2DqQopVtcDtjhUDJvfn/a
PAH3Fwo6Axtt7551uh3nY/ISR3vV/sndbL8+Z3W/Sgfg0e+2JlN+7vLXgw6k3PSCQDMxiV1vzrzF
ntmtECDqmL8AT6k6pIxBk3da2r+sPWwWtQlOzHIn7lgTe17uD25dZayotFaWGeDnDuIXy/vD7dzL
suLyq0GDuIqUlLgPpiizZWrBo6JRxnyAkGXTi5436ipeJhUUisvHBE3JyTUGas2hlCfa2I64KoBW
uA91pYUEiHBvhFt6zPKXMoMh5gCUEuCsgqbhgC6X7gw/tOVJKNdtiFcqQkiS9IxM1ZKuxNB9NiKb
yzAPv7tWJDyK86FqMdw87U+MrlcXhr1lo1KjkMFH9OHabJF8Hi+ZaXmv0aIZ0btk8Hvrh+Em6O4U
l24gewqkQErsMQLt3cdxW2U4+l3XwmVZ9re4WuKxPJdjac3nS+9Vncv9mITXRq2/v6G1mCGuMqpu
F686Ls39FqO2PlmR/IB93546MgTCAuvmjKgw6YLPJkCo4U4Vt8hHlN7441AoSEyUGP6ztqQkXY/H
X4RkCAOJ8vrWJ8CuoGKTvoI8NU3AfRLv+//qm6ls6IWBH6dKWLLtqbU15o99Hyi83GUnKvvDdARu
1R9geqTrUiOUpbKYP8GgwZvonXAFMnFUW9R7u7UpF0Ry13ehQZo1kxTOkyrD8P+KWc3luVQBEM9w
aVN7aMwuB23S11IGZPMOjkfpqTvrOg7G/BNDweGczM/rze6USdmTXp6xKa4dGC3WmCW1BJbfXAsA
nrcTXd+EofHmKEtRPa4kiOYU9V5zXBQ6Mko9cHalt0gpNEM1vp/BNLglmfFEvB7AxVhU20fjrLtg
iG8mW1yLjcq95wYd+uLoOcZ/qiy4kZGv+nBjLjVLBZbOvj/ucW/SUPcjlZqn0U90cUuArCNNigPw
f9Uw/Fux3Ix/7WAgThiRNzHi191OkQCL/I80cgMQSO2KIQt66zIyXXJ1+tHEbfK4Iv+N5q/t9DuV
vQzOzhO+R65LkI6c1GijFH0CrErBMUlyhxX1KnJGECZa7JT9ooMF1EJF3xk3N+LsKB58GimCk/++
orMOxpenpTGPx7gI6mv1WkP0M7D9yBY+SwR00szZuCcUplkLx1y+ryvTwiBFOxyPj77JzABaNd9l
OaKaWeaxwx7EGXMoFHKeKqgcunVyXYkaLrs90qyflCiyReUDbf3c2vJugarD1c2EQFSBhzF1FfVg
GfU8/BdIKYMwcV/pzdiqZ6vf9RwF6HI6sX/2RgFyv43XkCe3XmJNgJ9wqxFsCY+honmpGzbvP7cJ
GXfr3mw1/8mMHLWL4Ha4EE9q8PWEh/YUcqpn8OVXz2rAo/FWsQAW5HQ7NgZpL7A6e1V2YqgFy5nT
fsYY2tmvjO0aSbNgQjWUo0lIRmoJGTMeZCU+1GnN2klIuwUvoHhwnnkjh31qUhh3pD+lT2dYV7S4
pc8Lr2hVevDSNWZOzu70L+YiFOYjEVV0RSJZDM7xWDUUj8RG8w1VdNqK2ssLlM++jlaglCds8r80
igx2BlfS7QABnsX8OBbrAbkIAUVPd369g4cDckZxlPDwVbu/8TKXUwUopw/3ZSRq4y8icyT+kk5q
TlZYQ72Xz8Bky3hqJDkeJHRgTsdbqfMmFZenmXLsXgFh965qoe8WZPtb6ReKrCJkjhz9lLfnKbMS
fnSGjdOf5zDzRvS1lvrm+E3JDHhgi1AZoM6A9j9eurWst/A/w5FBMq9O2QMMSdG79m9fQxn7bLWK
OTIzujPY8KxW3EWvUICj5TeXPup+raofP8ceAvj9Oiw37jIwP0P8pFy3sLFRcnVihsuZtkYwYHMd
+rqnsVFugTc1UPgJMFY+kyaGowvPzg+tSvRua8AJiXCYn/1meqH2hBHJ5b4kFYQxRzIhe+PZhb7t
t+oAiIVJY9CdBi9GD7Em0o2QyC0BXUT8ViD4N2Q1gx6zaqybrmKohYy+1+tsSmqot3B0fBfyf9zQ
uyfcSS4nnxmgGSpelWvxcW1kVsd4R8uUI8OAi62WmAB9+R3UE21py5QUrmuv0187GSTrgnoENpVK
MLlfjWx4JUbmq2r3lYy6Ldg3MmqRQ9jeCt7twKa5hNL6A4gI/km5tK1xLcw2f1SMXYevst/YJ+KA
RxJHzxl3v/LKdkFIAhrqj4MtWewQu20CaAGhMpv6jr7/llxDArOMkD47F+RrmRdHCX+Xu9suZfMQ
NfEqt2aF11akJex+zMwCnqs4Dg/0M//dpshOpwKV0ASha3CJ/FE9b0tHKqhIgr0GrSGrjD/As0sX
iZpQ0meVstZJGwQzjbNHJoEKXccxggLBcK/gq3FKC8JKpBHUN6Gf+cf0zkK/wTl+Yh2l3HAG4aXC
pA+n2sZOVig4bqHa9DOqR0gFghb7h9rr2FGjySACHjLxMIUc5Z+iv5xWlOtvEvf4rGuVIRxjp2fo
cmrfU1/Njz2SFi4JAuiNuPelpEiNUcRx/LJze3+2u2fZ2g0USGjsuJaOcKuJ+M65TheOO4wJj0NZ
M9JV5K1FOJXUF7Gl5UxQmDvvU6axJBi007dWFeHu/zmAJ/vCrhDE3ysQ9MYfa8Z+cL1WcJ5mS+rE
0QAGdMVP/06yV+RX/6FhcdiZiosF7TCmcX1I34Ept7cmH9nlZJIAcOxp6ue6jNKKIkgcjCwVcK6i
9r4uSlRvF7sBn9mDNDtj7SBAVmitS9wOkSAr6ZH/WIfLV3VJo5nsfcCKZjQa6STEgRYcHrYbWvYl
kbgAqx2wBfk4V9iprYF6etNgq50+e3fRs2VTIjeKIZ+vHs2U8R37PcKDHiWHPx0uthxrfjbZX6Ae
XJpJZFz1YFqRAsGrqYbxEtkzDn01pUSiLGOm08hbP75SUPizfQhvoCEiRzLQRenqA3HQfgkAksAQ
RzCsKsAAO/hjq42k5Qa3irj/6HVAFqxJ+7BaoUPegjRz+ZB+Tl5+wYlhZw4Nfew37e0E4tuKTalU
hX+XZrnTDp216JtgTERuXr/zakTYVNpRd0hVmCXmugeDOxSpCdeEts9Q+Lt3IGznp5kZiFl/QHcz
xS5Tca+dmT+oaYJUnFNbHlsWZ+VmXYMRtPMQmkEnvlnLp/7KBqs0OzVwQYNxn7n+K/PAm4j1gmaG
LuQwcOm3Lv5aoOAdW1ltU6UY/+Mbx2vEYBA67Y5tuCyB5p6Y6ojvfrorlM/hzY2y4gq1LXRVDen6
BMUH439vXm+e0TVzr+vrDEdKnYuCf2n2gEoz1XoLLJCcB7xc5M2FByLX6e9UN4EqOr0fPlsmFPD5
8onrrL1O+NOLBmFV05DY/sgmPSV/I0rl+sSafSkhVg+K1Ij8mxgkE82UL6sx9ktc7KOx4Nx9ouIm
7tskt0DibzSWQdXC4SHlrsdn8omTgDoVjR04uSYR07MtISAqt3CV7cg7ub8mWWqp9AEs1Niwv1CO
s/3azn1C5pJ9fvz1dDYF6Kn6A8btFC9RHKG4PQkGBFzHSiiAMAaME6XujeREBzxkDOdotejqMlyI
Oet2x/NC2FSBVNebe0wluoTtBMxl9QpLxEBK63m3Nsx8klo4vnDFToC9iQMkKc7YxwY+JsXo5mmA
VubAgt5IB11IeUcip4tM5VTM+Pnm3iJVfnFTGG8d9sFsZHyX6oGBUSV1Hx89+23k3kpzcQKf2g9b
g3MOV4dVbnHkNGnBKuK33jehGrO5U5Co3s3S/slxTQloNuwn82LZKd0CNpjFopIeVggoYnr0j7n0
EDCw782PiQ103a13E0GQ2wN8mfuifWZvuvNrxp1KPh/KMO00U1m82/lNH0uWdrRZAo0jnqPrkLUS
A+plkFDcw+9UeoR353cJhx/Nnpcuj+AstiFx75PqDK+xKo4zxuRHFYWWa8PxG5rqpceUmG3gsoT9
Mw0+2IKdjsuxTYH0BnEw/sA7My2oGzkKI6C9t0JU7qGlmC1wkY9WFuIIE25rH9EHzDV6gA2U40zp
oRmqhfp6ng/8vP/0QSRbtB05yqKBXiGoXVE7sfATunumQIOJ3ywyxwB7UNWQRq3YxjEPcBfMx+vK
ko96CRYlSBD/zcPv+AY1LMNiN4tvyvB44cUoL3sycmFvmm42hW3uTgGoVcLQGE2EDKVTzKr2qw8p
YxwpZY2BTvVuKz/UigL8n0okYfz4U6tKsVqI+PjkyWikwvxOIRhi0F7eR3foWH/LKg46+hcDO64r
M7EgqAfmB8o0R57hNnLxHSmJFqjM/6X5Cj9FY9tKTvDNtukmnh8B/qFDDtGeVJ2YVVS7lu45ixe9
UWB7NzR9FwX6pjAuh4l4sgXiNdMetAdgiLNUK16Xl/Oy6Vnc2uN3p3ueG648dT9RTb5YoqZZR3z/
hRJ3t61k86LZLJnSXZPLwOaTyYFyGg7kqlm/4o4GgEtVAZM6ykxMtbM4G6wiowKqopzliDSKe50h
M7Uqbk2xtA31C90yroZ8gEHs6bbOyGKj5X2Loss2LhqESa5eAEv0JM2+kSabQpfwaFEz54CKVA2M
lIVpkqt/qq+tzhvq4XPO8/uD8U6BFd5pBdGCJaGG5OR9/TppC9JlsAiP7fE7sMBlmFojBqGr0Zem
esIC5tmYB9ysR2eXRuGHidH8gg1yJ++cGEuDS9hjcvqsnJu29aiHoXT2RQunBhI0P2bgmKw3eD9j
fGU7jMvzKZW9uZvfBb4zv1xHjEh12DvMaEoo+1uDSZJBWJnxtRFAtPVjw8jxWFsOmUIQe6l+qyUo
S4DR1pqnzKvmFKAYpV77rt1/Qy9eoB5fMqHBQ4A1r4Jsm91309AmeW17A+nay4ugUXhwmnWHNeJU
cB7vFprqlpHqYeI5nymqrxPKwSCaW+E25fiX6hOrIOeH+3C5ToPH9WDxtpfXE5bNtaFjlp8TkF8s
48eiDJYktr5YG7drXhya/jtGUgBy9LxtC9QFGR2v0GKvQFXNr4yMdRpLawQn49vTFUYmL8peZwln
CFWC8FrPWYeEX0D1XXp73l2rc5AJdodfKHgvWQIB3CUH92ewZbwUxTQgyQr9tTkZ7el+TRQrgzKu
ZopaTPUNAUM1U9bfErBNm+BM5T7souz9WL14kJ6hIbEPTpSYEFNbRB/RatlbDMVZ+aWIMxpUcVPG
UTA5Hq+uhQ3BrRlJWcxW+YRlFAka/sFO7bVkYHgKWX7cB9nj5OKKr7i+Ul08Na9BzM/LuXNQd0cf
jqJBvNg2zEBdeLUJqU1l1Dto1ys7+9XdvdithXQi6z6s+OKvkKgZ3RJsmx4c6XCIgZYQHoAn+lMp
1Wh7I9jcNcnRl+2610XevCYOQ/lIjj79tMvZVPWtE6cMx8OiISXc9V2wOVqFEXiLZDZMAGZOR7fL
0vip07W9iLt0ww0lIVTwHpGIpOrFgJa9TRNiePigddrj11DOvcpDtcwmv8sKgHbBIEAzXftOKeXE
J3gL4i1O7JroTtD9+kAj+JHTEV07+D+p/2D2PAAeGeW2/lpl72EjwWwWhIXlZjLYrXnzhRKtVzmC
1NrgDQiC434yBgHLg2GQbzONTTcZzIfACM0G1HKcCAPwt2TKl5SlVOjYhWwnnrPZ9K4vfcM9E5su
2NJCj4/26FTAVi70QgLEpf3K1tV+VSLz/1JKIoruOvID3vQALrQrM8Wjrh7D+OdAiCFW45Bw02AM
YtjjnMRnkKvEM1XSmCfaBpPvxHbHVK5BHLtRrR573zKKbZO2MD7dzcOnV3DifzgP6VWrYHOgpbCX
VLfAiXhBcTCMYrTGt3uxb37jmJo/fN8w1DAxuUlTojM4OGriuErlQDq9iZGAVOlwaVD+vo4biefV
uHSCrdMFpmSFNyoMrYbCliBysTQc/GZCEGadirTRxD5bTxdgEPI8GQ8R1FVDoRn3vJLs4TQ5VKqa
Md85mVz79qMsgoDFZTkzSJvBuKEHCRjkX84KhHw8WEd/vspwAlfXR7Oir5txcfz5yKHRZpDEcBaJ
60YcRaq+jHl0m86DMwmIxW75fYTzmE9RGhIqsd2vBOzagHt5+mVDKhsuxA7s2R7Otj/VUQKwMWlS
YCL6Zo0NkRLQDZ4ce1zrhp3pSiwOL4/Zgj9fLIoCyO8pUHzaxIEs4486WgH2WRr/15+4IGWbZ0Vc
zSNRdWGqE78rPasJhCweB3lRddwEt+R7Spay2+n43B/f456CYPD007e6IrHcQhObEDW4QnrM2y7N
pCLgCiC5nXqAIBs0kATuUuqM9ov+SVF34vBwRjeDx7fxKwzDbxdP1flET3HDlVH/eTwAeKrgzk9y
orc2A///GfeWq/jrdAr2Kt+ECmkY1Y8esa+NwHZxHlJlseaDWrn6z+ibZrIIAzaYkcXMQ16UvJ+T
Ep9fSTlGQV4LYpwaFESMFJejQpRDKoXdf+kKpNnXiNAeA6RHun+OWoNynfrRBLrWoB47WWZ/V9i0
X35bXPgcuRivrnO+FihM0ZaLDn16Z5YlhzipES8P0UxUJcIvABENUKNoo51cfP0g32B04x3LNqn+
6m0CyI0N5HcNdfhZvAJvacgLqSZUmepiAoKc3avqqa+tCSJsHy+Jibbhxajm3Ze2rolmTLFyWvfe
XFJf8XBevbXMIOP/ZzSdyLqNB5TEhtK4LztnlSxWQVy1uXSEM7bOfhfHeXsK2TehALMSJ/0APuo9
MEvQD/g6oaALIMAdiZKSJU2Vwlyu+gw/oIHc04dzSNrEUWhAignYVM75KN1BF8BdXTMhtWOzdOZH
5UcJ9od+w/yZcHWiK6/7lP0fv5AnfqOMZ2vMmMTjz/t0bWIh1dfLlq91BT4nPlhk7NlQ+/Dpgxk+
B53bJyES3IkeHZlKT9Pztk22ZVe268Q9XGAzN7g62zliUb48fUdIeH+3CTrUkOo+86R2NXCgl9Co
Ac1d33K/T0Jq94xKum7Bo51Hs7AGtWMLgdFxV8nXH9irT4ESGQD4j5jEXg+ZDx20W5ta0/6cvnyW
+FpCi8eja/8zODkCHEcdJ0I6J7cC+TMigCYlwcGnsKneda8ajQc+sJgQZ3IC0rkYtUJDr18JxyOS
elhWR/n3fZpuFsq0PgA3t0KPlj1cWZvwRsJffebTDWJpMb1SgWlg1Fn5vIgmXg+VBuWVk4iliHpW
aEAsgLKFoWWOjYh5rTh91W155w08iBypyw5EQjVXdIJK1IpD2YxB52A203LOsVOBQfcSLuGezUcq
sbcmgthQZftF6ZVw1JqzqB25XansL6lZN+KjgcZFhM9Tx4cXnj1hObMg1X6GkJWxcQj5ekiViNtC
xageNd5ETOqy6M3de93BDAu6cPU/mM+F7usaUJfuUYqlfttACyXlb8bsHbH2ESpm7vurQpXIpttJ
sEahJN+BMjFd7QA9XuC0KitFpB5GxrFgwlb6uLYQsrNA/i7lJsci+7w1o5tkICNFyPgQB4EUlrlW
N26L+nzmIWUgLHGqC1epQoMBObpQl00VJ0cCry5C4vo1SLeS+4bN34wK8AkxLAYBLRnW9yMR+vPg
xkm8XSp/6dI/g0asj/PYyPjzpZfusJ5Te5sWBNax32ATaTf7FYCzBTisPx2SkSxxQHn6u/toO8YT
4sCxOM+ruHHft2jajm4xljade5eeFSwjB35yyQ/yG99PRhzeLCfyX4e1cMUs5JSSEC0ejame9p+u
HZrqgRHrg8s53BsB6yB1abJCTYg0Sv0PNNVI1G2tvstxafZrWuMpSUEAUSM2lDHQ3rHKp+KSRksS
hklvjmxNVT9jsTeEHifgaCf+l5l7zFf33U8EOgXs9uO+MPeTwVjbQyRnIv91a8YCzn2hy9FdtLtP
UQ5V052IdyrC0xCSzfZoSNgGtodFAatBvUYrYO/uyJ6GZepodzr3QIoaAnVILqM3d3R3KK1OksLe
xcVVBW64hyIoVDTEJTVBDtX8CwYh4uyBztpkFXFfNeXQTzHTqyjzDLRYo6u1WAeb5RALbDP2WEt2
G+d4JPZJjuEew0upyZ7JVcNJOskO3Z6/15hlMZ8Z5WoV5MjQk3c9fpoYFp8NGSv31lkhihdM7jOE
aPGjVPiepyz98a9SKGWAC/6e49pCCrzyH1HJ2rdYJxOH/1qqXYsbHLbipiE2ieiaNKtiIHKk34hp
+sIrt2Y6CH+241xyfE2cfKaA0r6+JDHAfXeSr9aCLKHFJeJuv+J5S0vSak4gD0suLV0mAQFEbr+u
8IN4nTwkocvAcoUTF74gwKQktOvoZBHq/DWmisnN3rLOExsvtBQrV2+x5vQ/yomZOnJ8rUg3HAHq
otrjpj+H+4kGD+6OY0knALXHUljSAJUUsIAYb3p1eX4kt4UanLiXyFE17xCiGedsAG6OmLTWY35a
eYMT5VWWgMVKywGDhBGuOF3V9m6kBrGaiEMycF8OgQNm/SKQvPkjmqSDz+EwR6zt2unzpVic80Wl
jy3/Y5gjz/3tjxQMoADccTamjyh8EAnlvlbObQ2vGkILx5RFWhY0P6aXK0SfKKlPdtCecC1hPeSw
VdXZombIzAm4cAUe1RnOkpcmiBegPTH9nQ6dqVF19ktNnPV6er8FrguvT6oIRP50ivK0LbXWWq3n
Ob161aWBJoBWOea/HM35lB49Wp6ojg4F4oyhqRT7tDYRkoTTeB9JQOk6qnE/AYkFESXwvoez86j/
J20JIyZvmpYGjr3CCAhhf+fFKUDYmIjwoiyHBTtFI3DpfwHsqKCSrq5SQXMjTdmYhhWmNHZ3gBWm
pReFOR3hsk27U+gsModavRNQgqtz+QctTYT783CJ1Z6c0QuCfGh+vTO6WoDD+LLrNfy0ovu0+Ps4
bOg7x1CXFlsGG2pcWY4RNhXBxaQDEEiyQ1oevAy7u2LN2O2mh9wWuHZuSbX3w2lLHaAH3ZnVxvZh
GgEHhqu6oivNZ4r7JDyglcWYHiT3CSqhHWFAG9vpnCDz1LUmh0wNzA2QJRguTPOQiQEu43pcIWzg
UrRdDhYRPfaq9I8PniMB8y2VhlAptsLJBRDpsbmgbJSMcJMmskHAqcA9V7iEabQsZETez1BCgzoX
mVw69fnD2aGoEGNCTJONlfLquDVUA6vEo/Du2D+dOkDIOdgUrvW4z8VfF6nwi7UhxwrOP8Xip4gJ
w6oKGBL9ADPE41pWxMl6NntTgs6k8/nWi3G3ZK/Km1ih8AlllhkqKshxCAYZ5W0OU5b6Ha4IsH+t
/2X/shyqbpWuj32GGzMfqFCA+rLkNPMOvjfX9wgjRtfxhMlg+CCd3gAG5LVQSop4YmLAkRrZnL/4
2oPlDp8Gl4QfULm2XmEy6gNV5713BGuI3Mu2isqn06yEHDdL0RqDiiYPL8pxKpuj5W1eGeTm4EBk
rD9fAwRoP/ZITmJy+owXfpEVSPiD23HxhOz06J0ykdoah27Y+bjgPHM1EZQT7cv82KZC+mDvQUoC
NilslM3zrpV0+EFDsxasMOJufCtiEbtVBfNnMHc9hdPsNEyxLeHuY+U87Grdu/EiMklBa/95zEIK
sLKEWBakwvBdQm9PjK/HWnVBjPRZX96g4SNX5dfi7cDR98KQVzzIqtLmO0PNI3dRahNo75/gQT4L
Ax2oURtK/6w2Nz4cpwPMHYaG2MHuvHU8iDWXu17q7xgbI8sPEwqtn/nmURscbFEIOzt+5E93nJy6
9XHBxLW8LbMk2QDx5L+SzBa7QcxISjxEXArpLGucUIfDbpuyLkqXY3U7IhC2biitqII8OjkfUIKd
G+/omGfQQtLcjM9uQKxNPa77axofHv7luV+AOr38wGB2Fid5GhCTDgxcoHuXbBzw7MhBVUYX/bWX
gasN4ChJ5g37JrAZbNDC1P34WO9HIU7Gmnqd8Djk4aHMWc6bMKzlYFDSF6DcOpU7bZz+aGlVMB17
uqhzcOTo36REuDHzFdVuUJllnXcjWBFC/ROVNl64AG2uxQp2eB+DPYI9k5DGYY8B+mQ8ZyGe4ZGp
nzfjQ7XG2cqztaNxpJCLW2TdEY9Oc/fyFgX783jw/4OZa4F2Nsp1dkabstUtutJDGzgodpHA/eQi
FpzWgVCywwdf2bOrvW0eEFZ7SUChVdIr6zG18B6FYNLM0P+d0HyaW3dMyxhu3b0bjWQNmI18+rzi
LglQRwPumCPUIURi32H3KhUO2sDBcdY9sqSQ5LS7P/dfCNx5hupV6rlDJ+gfWehpCyuSkGwn4hf9
cGpPR5WrVbPPvOKtEJ+WGi0xoj0ThwKFlOWsiJvAgSc2caM0d/Qgz9fYxp5cB+4EHmTc61bLkoX5
gxT2LV8uU5I1AcshgvsUWdiV8sOyc7/kkKB53U6H+Wkm/71Neqk2Vh3bUYq3Fj8NIVWKmuVessOs
LqP9Cvqiquzv0S69zMZfzTe/pHc6HPN/vYQLJFbNqiDW2+InCz4lIZ+jtmXwBct2LCRRs9908/3E
2uLhTKL++dTLHRoJi3HJG/XMsylo/KuJJfmg5Z+k//qFGv28dJWypZTCojnTqmX0iB58FEryhQyL
WLgICJ8tCPPBFBy6oezEDZSNzLUYEj1NpX6pUDgaUqId1UJ+cF44qTTqQvADIbBgP+6iqCsDowcE
nzptjWN/g5BeitkhP4y0AJG7t8bjT9L233FGkxTlH+3dQcblZrQ82BX+A2+kCpAVvjf1+m3yeACQ
gM4MxriNIat0qxFKzCLz7fd3NBKJIhWkYPsc8EBZbHtUSVCCsB1qUoZleWlUVIx4xGeV09VogQ+1
HDWaTuipuV5404yZW3coC9ZbGAt9KA9YX/CUAos/gxu50cgbh992L9rpg3GROoNxXO9QwgIVmFdy
9pPdy6Kwy4BPZhs+FO33dIlVqM7ElIaYsqnHBgWvRR6SJnNcCAvMMOGjxxmkcZNuvKcJnT4RfjA5
mhRJsoXMPcgPGm4hu9pPZ2zdObbvJSo7zCwtBp2767X1RKB6K0xLDUTMQjseVgWWPS/JoTPpTWmJ
3sYarmWnlLfSWbKpIyuwgExHALzRRze9sBpjBBLdpSUemoFxBUT5VbRXlrdHjYaS7R3B5sNycZa3
VBNmXp0GNnNdmOhamJFKdmb14nym1jUga7E6btuxZhKaY2NLMM5XebP0EhCsE5IYC5HCLlDoYMYs
sN58rPsB3PncUuN4b/MIYMAEXV7x/b1J/2sx7VltNq6EDRSq9XgTGXMJEZR+r0zWqKRUgldJVv79
jWSAY2vmBEpFrTVIgognJ3b9Vvey9XQnGXeorJiUKYVVHo0moEMFDOed9G3gVUix27xXYfZWCMid
1J6GHfiPoV1UU42IUOV9nkPUCYo4OT5/2XoEHB+28F40EY0mISKca3gUmf588AxoGk399wW2ENz8
PJE8ZlCZIwFiaOdYRxbLlZLCtUIxNvHWhGTTyEFJIfMea/Ch0m8SsC9mLTwXWmZtAETvxfRhfPSp
lcmjCiFfVoxZREzgo4yX3ci+Gp3iK7GZb6hKLsPCDPoJ/nopN/JiIHqrO6oAiiymWyZYONM4Bpch
9TDGQfMmwJEMD8Do9GXfoeUgSIub4mFCvizoSoohqEYHZ80u2sSG6vyD6I3KuWcEk2vB2uDj8KXp
6bPOA/wACTl93UbWokI2MrK9HWaiB3DVkMaPD4ldxxq15uqc02EBFY+prc5qMMOhda1rv+rIOgE/
lN0QZP82+gr34pzbVY4tEpsxzvuB5IdJSr8qWTvP7zsXkLfoz/uGWDQO35U4SjMPwpSeT3/Tp2F7
JnLkl+dz4/RG9o3GEJLq8qiAPbYw6l6i5be2vf/So3zeCKpO/Qoh0jtqmwW76bZpo0bKEWOc+gDB
nA+kTWjRvWE7ODz/IvVGu/6oAkG0i8H+J+5RsoFj3UhGiuicl7lzAjrWPzXsxevcufvuLDH+7Go6
ZBWJhsP7277mzNxxPhhSVyiohNofxgLBG2c6i8LcLXKZRaswysJyuccLp7bVQf1bzLBy8E4jkJfB
ZF+MtBaLaq1w3V5HghEgOCc3iDZN5ZZuJ1D+Nyq4Qfv6YiQ9CQB9mRCzenMBwuMJpJRg17o9ctNl
in+OVu8VVfHyUf6VGclYHzPzcNa/b2Kml7n76ta31omKkTEx0DzRv/B88dFEWQtE+vERa8LgqoVW
ESSp6ZLhtSHkB+u02ynIsK/tVIWa3MZ251UQgQa1pgXYeHIh74lDlMBvgW9enxENxn6e+WWdItGX
zCxQBNVJAh29odziPGeULDi5qRyliKEW0DGxVvKs8iuY+dcd+/spMFZ/+IbDm4or9xBlZ+qhtwZe
Ojucp2nIof+glKPx2sqVSxuyfMcByRR1UMywGU4FVLm5V0kpK+ClU9z9/6EDrlm2J51vUdL2G5Ox
flL0DUzkVkiRfpLyP0E6TjXjnbMd75WjUYPIblWUNapnPQvxlEJ7ldWupAoY8pNTbsdSFbN551yO
EZ7lTXtisIQ8uewlKT8aB8Xs1dcxDd4gk9m5HClyza4sU5GFT+YZZ9QCBg0T6qwS2CcVpvKYv9Yj
DeUCccAkZUIQAY4n2DtOwgyTH570F7YFQuqSBB3VgkXDCRCEqd8t9H3vfRJX27omuISPMAViKJPh
qxa1iFxvgi3SGtzuESKvqzSi9qt3upzQjzFW2IE3TTz6WA5TFCF8F7RgkiWjs1O6izsHUaOgi3w5
LwlyryzgfnOgHOb4wyd6Z/gGrz5N5tbJO88lcF/oSGjN9J+n3qk2QxAAb/HGMX2djwlOkW+6jrbQ
y/PQ9GpY1AC5EI0tG/KDYXRBk48jUsHDkiZK38nLUWdyD/9hXQeav3rYBnxW8gOxegurnElfOCYW
hBZT7ydH9AJxTriOCnhS+3xZ3NfnLd+w4ywuh7hqVm7B6tLyICk1l9VCQ2p6vzj1c0quWn8BfZWH
TybJ7A4Hj/sSHcEMywhd3k/Pg/ECbXRmj0BXYq4C70BnYceAW6jnVaBwaFMLouxldPq6c1YsqwNE
DhK/E77USIavTQBMLDmHYvc6fiYLZmUiQyToVyat16iAqNJL/Y/Y/KOjVDTLq8gbeKoU3QibnfiJ
RBJYeAXPQ+7MzSZ7no/4n1gK3Fx3fYSDhrJhc1L1VKYclG63A5reQ9Z4273cfxFBoYyISIC5ycIp
l6zTgo99jsHvFqoouBjs6zVzv6kAyqedeOmSyS8cI6CQ1MPIWCGWuu1REmdEr5+Ivz7ho7mMuq6T
j16E5ELNHk2LVMkmyzzADALBzPfd6iPudsmbnScKSqd2foQiXMb3QQ8QG2lFrWbkj5YKu7Bb7gvY
yDA0OY+cMxF+dzulXiLHq65AI6Gy1eRvU4FnLOO8D3BxEtwFRtMZhNFUYQwgxeETRpY1dLG6Um+Y
lWsFhszLwM5avdmlF2quOcgG3pBadBGhWfASSyoKya4KhJICSdY8f7gqapEuAP05e+Vd+kKJgXLA
ckZMcgwWFwuMAUaXbFI3RcbEgJHNYMc+PSAQXukLoPObeQsfq6l8xgisxf98Ii6+czA5Cfaq3AuW
NWyk25FHixJLCcbBpi5wb4nBPSjQEcODolMhofD7SNHyR8Xi/hG2tZlUryblsBMADjWTqlZWXnuo
TZho4CNlQUGEH1iTCUn+pPPNlfGVZ6Z8mY5SN81x4jdS45GL+JAAVVsnEqRfHkoK21oTO+ieWYaZ
JHSoaD0h7bh2pMAH0s8gTR8sbyhUajfb47jRXHG7C3iinQRAtRa43phaDksMSQoKtRqQgPXO3LUz
9Q6+z2+8SJ38Lxs0Moi835TmxL9UVaxEIbY22lZerbZLxf4UW6D5sk50P5+tfWElcLc9Ql+DbHui
hElYV3Q+XOozQ6oZsiYrgodbkW4WV9ByMAeTJijyGioTc1M/M0yhJEnnBWXdNPTIPQLEJhNfvb1d
xtTazVZE1/znSIOiTRATM/D3Nh8I8dtze2SNjV3U/xH6+2F4X6WlpabTfNoCK2iBSowq0iQ59gWT
DfLwGUzeyjmfD4H0uSiFyFUeCZbEmf9WMdzaQJejUSWOaOZQgWlKl1WLOJAzgMfBFARlKKO2MQVK
M2QnqR4enxhYE6mwnVU17aE+UbBdZ59RePOjwySBA70bSicHDHlfhQJ7dxtohbCDjzVS3kQmSfsp
h47FWYv7aHWXuNmOIlD6lcUlaoxlZczGSUey8h+4eEIDqT/0ZG/CLF0vhrj0y0SPx1umLdGcPUy8
TZ3qg7MsS/nbY8ZcRTpdyLUbH5T0rptSziiM/h+ps/KvJZQlApc0L4eRkLml9qYixsByE6zOp1By
2oYfSaqAAWvCpkwa3LCEWl7IUAWWHaFTwYC5eULMVQ8WSBXalZdR8e1nKJQMhmwffxEnpU51yHy3
LaTgrWWX51FvfaE6+gXI31B1V8euzBrZV+gWr2wRVPcmLOZm5p4YTVUcbZ2FQtITl6PJna/ailoo
6A9PlbHPsHa51qQcz6AxEm7we2v+Lq8UrKztu4zWf2w5CpGw2KH6dBFyh2zmShySgCJ1MXicRmR4
+u0yK/ivlQQ+f+RRWrl2ZfF4gIr4nwbbeboIFd2SVmil+ow2efyRDwYbwZhAi4VUo7eGUfZg3NMv
vCBeXzUaeFYccIyQUAUf23Uut0DBLvBnszzRWaEiMVySMqS+hmJyhr8IlasZShqS3KBZtxB1g7/A
GfQkIo//BLwFcJlLufeCKcDZaSrSJ6w6d6JX+sc2o67zk+UGyByvHwJR2G2h6w8uWP+NA2elllUz
qzrmxxjCgXpF7LGBWHY/4uTqToh68OHlA0z4vWbaXOHpZWosZtpNEiaVINEMYMjI8pC5ZPNzNYS9
YtKg5T0UB3lfv1qZwNRTao1J5YcmoE0p8uhHAEyzxB0m/LHvs+5zc7Xxudx1jYy2Z7QJbYtDtRVM
KIGVyVKj1gQ85RYgj+Fw/LBznzBp0nfU7ekyFivtIebZjvhHLnImnXBJ4uoz6aDrDkR0OLZqGwwX
wAWeLgSVHK9A8fKhehV3jEmLopiLOAV38jTH7D6OJ2vWDlt7g9sPKoksXL6ZXlAEu+5dJJuEdOuj
beRmvxE8M4+1rugPDQrZdpUup8MTxPEQUubzgdkeWZLFTUOee7CVZO0il1m245T+XstCPCO1hmoM
qCTKF7nVXADxfW1/Rh65qDhlIfrCCZH1bq1ypzBZ3+ERFPPBdHkxkup+HXIVLaVnCFGw70cjbGLX
HACOQ7IzNq3DFamPHB5NkpL3hWT8LWFOsdAj0kcDdy6qIVcY4zgHGIYpTrjfWnSlOhQ7IpWkNkLc
wpjBG5yG8eSXuHr2+aln1h1jIMEFXGkomcDH2euOjrsCThHwWl6QvxuFXRGP02JAYRc/iKeS902C
4m8yJDLtyOrg/kf4p2NXoy6NfwLK1FsTwpdshpNt7CnePuWeJIzcXpapPNcFQjExp4S57WX+c/lf
T8JINPBRbz23CuybHe2AqKIeM49q7rtQQ1sjMgmGz1c4DkHkB0NTuBjfQhaHifj84S88Oa8ECEtT
cOtxgOBlTgEDerRCtt0bSutUVBNByCrB+xwtvFdoKulxpnv1PnY6YonOiilX8xQiiHzlrLOQomxy
yXBltcm55c0/7Vh5UfAkTKoMo8h4oVCwriTMJcHwQ4HG/kI1Ao2k0ng/5Ti4Oq9U22XecYBXBwsG
I3G6TZyC9H1Zq99tmOM8/erTiR8/8+pAkSlIt3yQOeELHy3hv+zXbo0X2C3dIvlueQzVneg952sF
WTkLoq5cLDT8m4fATuxZoLZck2+TqgT82iAOTd0mZEL4u4Puux28W9cABtU/dTj/DoQ023Go0nMd
wvVQpJMYavqv3GeRcLXm8R0h+mk7ZoevTdg6GbfJeGId1VTaeyH3h4YfOd+a9tbBqXYpKkQZeTAh
7/xc4JfMHKadHewpgr7X58YWLS5uphmE1jFPyswyU52SX5wQdvzFBrGzbHQ6b+mBqSb4KH8BfG8Q
Vf/SIQHFQEbSt03pB1t0SsTr4fBzuk6OQXQofzAAUWxwraHpOP3mivzREao2qSTIXJUVM5yPIFjx
LqJolC2CmxBDRnmESv7n42kwbmpNthnWv+d9B0YLPtqVFC3Mp0TGAUp/t1VPs5nar1qDBCVvWQeR
cb/Y6MgBome6Xp/Q2k2h5WBVx5wUScwWF+iViEuCftdwiT/+p5p7tppWt0o/+q6P7HfTUo3v+YXC
yGzXOu1O+pyU20qzfytrE2g2xBwB38zVwecDZMSZKBGYiiFOOUNqIJf1jhtcQ8xMPgx8atIGgMFs
DHY5XodsPlxEiRzSPQwT9TB4dyMlH6LZ8GJCYo5puv+juY74irTa2yvKrtjZDTKyHLVIk4ciJeNv
wuy0FOguS2YThpK4OtnvUhXIydAnt4Ss62TJKBWkDMoP9H4seLEvkXlLWsdOWrsNB5ERsCK7BSBi
aPGkLV686JoJwCT81JP8v8R3A30lwq4DJJ2eu13ChoMWUDpcyDhoMIFAaH35dJxRbI56AivIAjSh
SRkg5MK8TLznQMVDlPva89A0r1nFhE1Fh26ijBS/dkV3KmpqRv1RGYmG7pQPiZOEwnoHvkoVEenL
p0M9v3F7AIxiHowcjOzSDdW7NaDy44pJEqbed2LFQVK15tfpKVz2Y5UsSvs4CwfeOv3LLdjukvrM
55JMZ/GiqZURsknW14WgWeG31H/m8+YbUyCoFegrPD19XBSdWzKVZBKCKCyMqfaBLc5Wgv1COlhm
56m9aUub6iirSD0AzGPGrNxO2cc1om1CJcXbHulw3GKB/y5KbahTayf1p+mjkoSTfJZZO3jotOao
Il4HzTEBvCjMBGFu4ESPJvfhp6CiZx79Cfr6kwLwW7xr6xEvCoZiZapFPe655yZszhm8r9s5PbuY
YQPpTO3s/qoqfze5ytpyNsbEumOmR9UW6WoctGIce3md78U5a/NsgKEOqWAuumWLnuD59h8gPqA7
ZlF6le+MqxYqZL96gJkrzIbEF5xDGHua7tE0z/InDs5BmHI0XiXE+dw5YtfdCt5up3om53qrta+J
cojMXD7j9C5Mx6CUtn/ND6hQ/xEmmn4mj68JNSa9UJ3t8AIHZDkK7+hMo2v5q2ldhx714y98znmv
96j2sFgdQAiZnYfNuCRdaXflC7el5ohUKQOxKpjaV2jrvr7taclxv+1xSKcoNqeAVDLyynVulchz
qgqrW79roEWdUzDUtISDaqXKBjS7TJQt0fplsG8mAiOkXS8CAVB/NPbUVXnSIyB/W+dO0akTL2lP
rQM7PHrRuNKke1oondR7fTQAJS4yEU6+qGr8nIzP4ehs4mvPM/AsBbumXwwNS/2C1LmF9Q1fz0u1
kEWBwW0v2tFpbYqs8YvDmxB4cizprpnnvycCiHU+zdZHgUznIG6o0juUzl59aIBPfEuxWNP+mB5p
Kx6zQ0x6YXXsSQzp7WO9l2AhSO9K79B32gDICnNfew5UQfrOVDJFZx3zfXdNwaF5qV2aOt2HgplP
C1MKaKS85wRQDcVj4gVWv+tv8eLXGupeshnMr38aK2127WyhiBwj1+D8xehqPgwc5jPvmTPJa1lT
Sa21S8yTfy7Qq5gIEA+KXVVuZ5qQAX9fWlP5JsE3tW4sNjUMKQhVsfauSwNCZc/C2/CT3xioxtBE
VsTGudBFj7NNyYskK5hMC9EiQIB9OcMCeGBkpVZNl5oX8//R/eNy75nctytMkbXVRYo958uGj6b1
Bx1vFbCJGaOL7HjnGbTSp2i0qomXwpwvsfg8oCulLhI4TKJTD331Gpi0p8/NVNn4UJs6HgwQGuw5
CLxI+NXDdSgvNowOKbFfUc8/ji68Hc5xNWi3S6CHomaY0kdN+ePF0ie619dxSXG0ptLuiNPQ0c9i
BXH2HrFLNLnLaGooK2noTL1RBHIELbj8Q7hkrk4ljv8WojpnAV1PMCqCzy+FfdRXU2NuLz3OIr5V
U95ruBhVlm7eIiGWWKNEl/E8NdrlG1P4MBhmRj9ASseestLRliKGsLV/J2AQs56xqfr/dzDX8fca
SGp6Tiem60kv8PM2JzdhzGx0gQwA7uQ13Thr49rGG/8TKrqB1a6xA7awdYj79QcrRmmz8VZ8bUJo
atZbU+8ag9qWOaW5SqoPP0ahz4ijPDWCciqxNH5Cdcoya63Ttw62Ofdk1Kbj6nP3JS1SCnxkLknt
wCNlp0i/YNUyR/MpIX4rcY9A/NrDpv7Muc6wZzCPPF+fmWo5Jvh7671Z8ffe53AxlrBd5hYAhFL9
tpdOb0eHN2IFuRdPiiakJBNw8ygoWHU+HcSSrpinDiAEYx788nyXaYdYUtrvQqlP+gJIzP4YOFiI
6WJ4yvK+SjGNKotLFgQt7F7BVHSUjuGHOpSmEmv+XyMlyvZ38ShDKWlSxyj1sU/3TlTkzM/nfx7C
3yWyWW7YmCpfzFUxCYUF2tsl5bV63WJffMYD+Ua6dw0fXKkHRJ5j+hXj216znPqaIDqj7mypuAwM
4HXTELLDEuGviXwIj8dI3vIe+hmQo9bUx71uz91+/Y/uAkEkCzRQ0vXWfpv6w422xDa9VJeUJgGS
TaLHaSzzey5KTfS0Ci1ZZPyfrevg8TbiEig9caM62ZouKM8EZ3N1H736DneJoZNTmCmKB9jk/dxR
RKx6mp2raotVhNEA+tzWkVfJfAjDoynMbGZ7n/4paZSc5oLErUHfGyBC9Ec5EoufJCapdoUEhyhh
scgspZrfQjD+A+YQ3vflvntHkJbHR1i+8gK3D0FRn+RdktU3WkhzCdGthaVoAWF3GQxs/R9eNGeE
sjpxrfqN3iPhgQg4IZrP60+5j37b1rehXyObiVEe/lEQZLoYDky8F1e4AwK18fWvpxDfzMRJLVxF
4QRmFOwvWn0n3StPy9WVohafctoNekvCkaDA1VJN+gFV7hVcBm5B3goFTXycFxaGm893wYTcoQgO
9m40rl4I1DoygVVy5mezXMFKlYXT+1Rj4a2bsh7kzr48OvpJaStyC8BfkrlXGTYqxcYCjs7RBb/F
IjUvNRUn8UQdcmSzhEdAarP8yxGOwJVtImRnXbzhbgkVaHpp9H4ME6JtUnA13w53wi+LcEMCvGXw
RtsiA5ioFn3/xr/Jq7G9tptgxsXMPSvVia46eOiJHB8BU4HnU8Q5+kLu0/0V1+8mcM2Lf1nyrHOB
tLkL6NFoqZcpTfdvFeubYYQSo73drRFAeeytHjMPWPFrbl5SmUjXIZXQ30isXkfIjJReJEWg07z7
dqtCPjgjypIsS70Jr/eX3wIneQcMad/K1grsaqy4O8HZzcwx4lER3HZw/5cUwMtnmLkEq8zn1Fjn
a56NSL/k7uPY/pfzzU+1ZcUrRNNkBPrUXnQ0PXvn/N8TfhjZpAXIritjJ4aU8vdJH2/JXlYqyVbn
0kp0Kq+AqEHoC2bIqYbjNqUPPSUDQe15jnjgtdWrn4VNq1Ig4NDAZAApGSahgNmH8Gm/WkvYR+Hc
iGJJ73Olyyz8XIQ/1i3Jo4fFw2nIrg+R+AzByiL8UpejHRpeWgaATKOaVoQUQxHyFaJ6t+fD24QI
1k4t6NcT6W01xwlsWr58IqQnUCHCrM50agkknhk/MaXFZUy++NxMYQqHAw6A6s4tFxGXBjuODMHq
4f6sSu7jyNAdywSQWcf9XYK2w+mqfdo7lqub/W3vcg/iqv+gkHrqbZTYLCfdQbr9wvK9P93UPn3X
+1GHA8qalUUC8uVC0aGD2dMxiY28NxXBXQlfbOk6cfNerUeXA9VcpBmUa1K03xzM876ukkJn/DVN
Gq7/fN885BzHMKfJEsDHjwR4Di3YoMBVoF/atwmMv2sNKzz4u/ISeWGHgYHJd77e5iTDtGg0SJPE
hiQUiOwo360+g7lXNMcqCMSiZ/AaEL98sso1BE687B6oQk716UP7Xl//uYCYXvVdSlh1RmPESHXX
H2vCXWdPcYIERAVcBF2Jf34b0f7UNE28evctyJ/QdfagaiswS3ct+lqEswt6ZIBzPhOnKHQVDPaH
oAo+30fn3WgUFeYFJ2OYLsliV7kPa2agjeu4qIZj6k5M6VzP2lnmLrDLxrPsJqGjUPDGTAXb7Idp
2Vuvcnk9bvJPr39Hc673dQAVXv7ibpBgInw/qD+tqFeWgcCrluOs0zL11w11FBApx3EhxxF2XwB9
+KFQKiGe8UoJfks8sLSrUvOzBlp0hkGnrnOSSkorkfYv712TKQ5s8+GwnLmOWEyIHOPTU0ZnX/Z5
R4+Ss+SUDc4rIVHzaQkDo6yE6wy3J74Dh5kGQSh5ThRhuwV4jnkW0Fl+k3zuUJkMWiG2T3qSFac2
cFlGSiNy3QV1w8z/1LSKwju+NAjb/Z9wHdmWKLgEVUGyEZDNeQ4l8yBFI18zf2FY1rQKNRJu1b4Y
wXSGvsAnXLkg3ZRbWc54OjlzBuIe/AtijlLvd9n6h1ZnjveVfRZMk/3LpOln+qv1pd+CwzAzh0Jw
NGSM94EV8NAXDX1PrroRlYxZZ3ZpZR3vZO5VQmUYJetr6jt7ARvUmcqVaGtHhHDAmxHwLvLYzt79
zu0uGWpEwQcEP+rJ0GDBG4v7qxkdEtMAYbCHfKuAFxcgJqGpRt/Nh0v0/SukRzW7rQAd5vJcX7NS
lYsKx3WNvFg3k1hh9bSGkzduIrhC+if9sI3ZHjIYrHBAX5CUhx445CKGWINfRBUIB5LtvjSgmRBf
3T2CN5SY4c5g5EadlUMlkFoEsN2hkaOeP8Xl9UBP/Ua1fpy8TI8Z5KdI3u9DHZtlBIs/QF0MZ9VB
3J5jyp+wBxPN+1gMFF3mK8LwFZhngRHk1tlcUDhEMT/5dm2ewgPGx+0CpfnjdIPgiFA+mwItBBTT
/qsfqqItg6Ex+f5RJ1EN0NzE3QN17SbR/i11uPBR1QNY8vy7MT0cf8grxTPUTGd/IC4clpFIAbkg
FPiCck7fm39xwNSwIvUMpjMdVC4GdpyBYnl/1oPr/IfrV2DvMm0KyBlY+yWD3GgIVHUWcVDfmu9M
kpoW3cEXC7ZbWlM9YtsJ4AigugYdRhgTc21lkqu7521TAqZJvCCypCLLQr8IPk0y4vdh3LEY4SmK
qw3MrgJn/4QeKAsyHdpM9zOE38OrVf348TyCaUZrOa38XVPsUwe7Em6rKBrphWNigy/ojmVJyPTH
jofgxwgrGfAc+py4V7RUC13eQeVSyVAxROFGjn/W7M79j4lpFT5TOWg7dWvKiuaWWi0YDmoZG3lr
mGE5HKRytXzWWC2PnQmRHhVXv1gI/GSsqm0F2ZVfeZCzu802Lx1bFPeovngsXiCnqVTmBk2EDxFL
ix2+yl4vdI1llM5bQV0sWlBSF+x3rZiWZY3MJFKRTxSdddbr667jC0D4RXQPxIc47MOc7yEk/9Am
NQUfvUeAoRq3hVekhMPMfKvWdGrJVczwmw7Zv0WtsltY15FboipIq03nSkjVN4Hus/oPk1hrawWx
mOcjrhQ4l8oVMssbI6loqObARn5CMTbj+dsw4rlf8CLzIvdcWxREx25WUFiPp7JKTosNpdsvrmkr
GeRhkUxunPa5vNQhZ7SnpP4Z2oi4hHS8zO69XuuEYokhGnu9IgtZ8zmVHF9uLYLxOU/JmR8ufz1Q
ZbkU9xLwwxqrFzwvGsh6B3IpRSpI3n2mDbxPgylAI4U6Vs+NQKmZGQnS2eMBbH/8TtTaE4ZDHC1T
W8HjgV5DbfOws5EIUWHZpRYq+r4JTBXmaYAWiLlOLrVb2dxfeBYn/r0psxsUDcYcSN498E/Fe8/o
T3v5jZRv/TfsXioisM7hLseoEBnlJncWSSOFNmdozY34mEwkrxt6em5j0IfC8FvLIT1fU9cc2nGC
YMYR553qnatsqK8WUpCw9c6KAzyVXjciEZDmVjVncUYj0Ahu156l0gLHZ/DNnmE+9oer9v9BMvfF
AkO8i/qm9WxSrY60ATa5HXLtHep9+7J8jhY+0ArxpgjgJfGOHy09wbIm1qmaG6KRtUvtO8CNaII0
kpBw1W9QDtyirKvNXAmjr+Tg5PKSsd5Ed/eCCryC846yOjDvkPzE0TevAt+JbI88Ejo/IElo0Qgs
l8ZB9NKSciIzanTqk+ofNnS0aw2gHr+WXWitcxslWPRBI/idtAzm4SHrtl4wNpKbs3gie3eOqZYR
pskkAZ3+SVS0dFR3P5+TknQOSNTfzECT/MGcaJln644PvtkYK8TG0fiF7Z4PonPdEM97as9JqGQ3
Q/xupGWyJBzBTw/vjMASAq96SzqSE01fKgur8ktO1UnpcWubL20IG3Vdd4oZEEWKEIewxp558lQW
WyQvZ2inGGLPRWq1m/S6vpfsmiY6H8/+FrBImitqMJrAW9QYnkBHkszofG89jd7mCHsaSBLq3LCJ
oGzAfqZNvYENJIsif9gU3bN0Crd3FGzruwOKLYAW7qwUgHebIcEidxRWB9J8UwqGOcB/iccm213v
yfE0WP+2cNzB5XcwTyqjNznd9u0CjfTO5lHkR8xSWR26Zi9Op1QKcPddnth+x4Jug0r6BLPkoPGW
1nhu+mKEUyWIKT56N050wdlxEVd5f2xlIgEGqAgidwii9uOmRsJ55KW5s97yZNkQ6S9bPuO14HHa
q1M/V1SFk3lsdg0jHO/XZqwl++dvdlWx4/e3c5kA8Nt7XS9sabGWcJI498zN/jEk0HuhBTcG01oO
w04eaqTDfbFOiPkcF2/rBc0o8VlyrR/nJkNT81ztDJSli1zI0uxMDPB9TlYYw6Ev8sWeM/VTiwDN
3QhsSqCCCrwhb0oIkg4oe1MpUIe+nQnMHrOUfc49RRrxMCxrY+BMyVY1F1SQW65oUP5e38EP6bTU
rtimXFACD/rsaFI+pV/zlmoETBMBkGHxWH6sq/g97/Aw91K2H14AzL9OHXLorj2VKIn21F+VDIC7
PAIx8dNXtRaUdlutIwDqOvhNoR/eEq1RZnmy82GEOvez2+0vqgE2qim0+GGs4WVMLMwuuMk8AkQ8
ieTQ+MQM9s9jwQnRK85usAAbC0EdWhhg+LHYl3tPDSjUaMo9ta68JVmuNtd8gZBEjHA7rs5j5VKg
RhgzOD32uQnUpOMpDWwqooEBliO/RliLOW168DqvEqcK2e+t2T4oC0wcGPCDPzZvsOhIm1uKFapf
flpJqzuLIg9r2/Yylj2bRUiHK133vFBm8kZ7DcQ5llkxxuMgRt/dOeew+fukKMDPyLJqz3J/RQ11
GXnrPF83ZcU+wVWawW7SiB6BEIuUG//rWxwchy3nszYS2t5dvnQ/DrQ/HoBgtbM+39FPpzFpIXcD
RGTgCUHnRWfMkn3KHV3x15PvPXgvgBT+sitIfT6ge1IT6p2RT0qjnvWdQyvdsZ5oowdby0QVe254
SYhwkSnUqqx1U7NI9ZP+ogGWYQOW+oME+K9iF3Hwb4TVwyyQVtwamSSKTWMy+DpQXhZ21o4dh/29
l4A+noyK8nBl5mbt1v0VlrmwIL8V+Sfy8xkxbOE9xVbOWX9/fpvRYnnxR5a3XNVNdEXMg2flBPmt
1wYDSQtPp93Y64FK8yTCxw9F+0s+O/PE9fr9cE+gVkcMADuypZSqsdle/QNF9IaGbvGbVhaBhh91
cZ1pNHAR+0euVxyPbdk0vbvzdDNfheaTm+9uMEAJe+9mZzLUsy40LFITZ+nRT1lSnhdDq5zrK/Kb
5kcFc2UWtbf15KsKgw4DqJvEBu0wio+Z6FvkPBWyMaGOAfI7HD1tz+78kCPMEA0nMZL+3Of65uvK
T9rhwIEk/A2N2wlMw16EXlCbMI4zLdimNAz9e4//l6FI8VndO/YRS9cYbyELdXYZgyDVPLzM4SH1
KTTFIuDI2nDSIbBiCWdOBcKiNTTUQZ4Sye2mVpN7mGtFm/HchXg0E120Z7k2V2H5C8/HlGmmDMb6
gzmF3CmArq4HRg1vEChuls9/KMns9RA6RSPKn7ca2msZT5pD8DxTEGG1QztuOeIqfEq79o2AQNnV
cDn9AlEh6wRcL2SclzI8VEA+ZgwiwvCXPQI+WB9+VFxTK3bB89r7PMFf8Fw4aNu3heB8qHZL/fKp
iW8GGQA80zaBycgzRbiESft3DNQnMroTndR55lvnT8ictT3AQYD+qH2J38lbykuqbH+I4eEupAjf
HK9nndLiZYEeS1snagptHBjeX27LREFB2Lv0xnhWBBBLeESdpgU8dd+TrRyrvm83+a9XWI3VPrqt
gz33chvrIIGQeM8GwjewUmLpSPy9LxQwJ6EKDn8GbYw0wl7b3b22PbdcW71447j0uWdR3gBVHmr5
E6oVFuOd8gZnZaWcBhLmJxwo+1WQOKEryqssZLWzHe16l7qhKIVWO17K+t1jsv1UvxAX62J0lJxU
bc239m2DMV/shrflq87KErsuVD7jWgq/tnflPJ8ZSmfEwhJGAq1JZ1vJnNqyhrhLFp3t8wz94Vj4
Dl9vqaLm10flH244xJvBYuvehSr/PIdH1nQe8fE5LihXHBO1IWJurQ4oM1DR86nkiE6zGB7sEc29
k0h+AP/HE/2uaZps6n0Jfr0U+bbzp5WZySSlopGmtlyKzTC/J1kGpK1G/A/mjQYaSCaLMvFzkgNM
FIHHMhKzqi03WOuG17WHfv2kHTsJL9QhEt8PYoIpBUKJ62+ruSx0ED8RkmOhEWd293gv+5zC+6V+
ar6yA6pLBZ3vEhMcZpWj0/jNhHNWHbAnVio5WqHIxd2tKep+maXfdKzrZc3GrRHGGsH6j+LDV63i
ZGOVlU9qn5ymRxdeQb1J6WElDED7tHWQ+xy35Rh3Q+k6aMhV80B75li3GmruhuwLmoihF+zcKM67
lwwts+MDevmHMArYwXldnYlF5RR3nqidoR5LWInUGw3Thcdpa0fGdq0e3Wj32+1X8V5D/rx2E4k8
1eCiKlJAsoE0wNSfhHjRMLdVCWVCtn+Oa8x8rn6l1DML5YUoYsnaX4TQkNjhZDU8Z72UdLXQj/9C
0zLYQbIr8TvVewMRhcYLGIF6vNjQX6mCXiIyMi6DZXqQF9r0GsGbrO+p40MF5VuDKk84EVcinoTI
dHutt2lqifmsoF6DOHdkEt5380yWOX+kA5HX9+ymnEHBujj1xX7+73eTTuXiRJ8h+mbSsvvfocQw
ActYY6VMxX5DaCpVk10/dmcRu6nnTScfEv5/Ek3NpJKamcsNnBqSe1OYn8IGioJG5oQ3pcenWMK2
+4+Ht80mg75NZSqg5LmyV7WRtyiJhhA8kYBc8unSfb4oAJwoOdLrRDUqNOx1yY06RYq12LR4JbmT
/Iia+Z8zCrHf4MWdrbrnHmHXR3XnTGO/AopRd4zbNrhlWqIhcpiCel6HLHf/COmZZpjyNqQnnvrn
LMp9t4C/pNHrSzUQ4S7A1Iz6WAX7M3SlWw8cj8wTP5iHkZMtNUQQdJ2BQhNI6eVTOFmfa5XMka7P
5DrwzAyihsmZVTlU1VwALPTL3bHIxDcPtI4+aUm0cGY2qY9W+v82mO10PIUxgRWMso58XUM058a3
0GRbHE8qRbAy757HFVYV6HogkYK60wr89csZtnzt2yIn9+uD+39bm2PvjP9N8voQP/RWVLNI0zme
7IwQKAiJQ2XFSFuOZDIJErUGj/tbDJl2Vte4JXSH7YuTWJ/eGlr0HNWKRvQ3YzhAIrK8REUonZAF
KG/5T/dVir1urrEgqJ7Ki4QnvLI3ieFD13VyXI2v8qpke4ppAOELDCb5GJuSIGbwKsR1jYk1YIfz
1/cNwtaepzIXBBVAv3TSBkWoVjM1+Hod5rqy16qc/lbRqoqiiNKTChwkWAn57xzjY86nWogD6osh
9pVFdbAWI7Xm//bcirPl1cx+OTji6TUg8mnR6+1VH+yL1frIavi/lGHIDq7eZ6l4tYiE5CiF47Ag
Ez8gfriJ/2RBP3lBGFpyrL2FbKpkejBOMdnaahEezeKlJbXxdRouC3mIPYhPVWowf+MRNwK4kCGG
M59IWP63zgt4V9AzhAAPLIZx7WQP9fQfINQCkbsEYwFEZqKCSunF2dlJ6ZF7Bt/mDjm6QQiViJnl
qstWS4O5kvoFtjhGvBwYx6iJz11+azUN33gw9NITr2VqCp+PFR94gV1hzitvIoLQ2Kmx9kXflpRx
E4VFI7MaSdDsUr4uNgxIxN9GRaRvJONZBP7MYdWDVrLAe73PjGfv3kYvaWn/BXxYi5jIzO3BtnY3
Rn54yMyhw+BrMDvj6uaUanVVMowR5Lox6xXmqX4zl6f0104GCAuv9LsbToYd2ssfBTNPpLyjiztQ
OVpyk24+zQc2R0bmnbHxaiW1SuC2x+7xfbMWoWf3tKLLEOsjFQ6dtjKyVwoOnzc3Ml0RSYmiLYhC
CTJE40zqeG59rvBNXajLksWA5twmTVyCbBkoN5p8uOd/IFLgAOmKrDntDzPu22rVmnr/HZp4PB9A
uCS5WeLrd1JiPkr0NPojvS5mKCnkUwTAVVO0TTCm01/1Gnlu+jOSCgyvxIN0wDnJtPkYzGOxybHJ
Q+Zl5JCY7qCPsF88vjeN/HvbZilnaH3kJKqGqeoUaJqcK6dk23MrejDdq9PcO5S52w8s5e/+tf2Q
jeyr1WmmVZp3wPfC3aUCwo0xz59f1otxXLlR1kFuGiXvSecHpLWgb9WwkPBYFegfn66R/K4NFYt5
7Ydl8fr+sQwgt/GubkOl8Ov2X/U97rbZOpQjMEGrypEUf1YxtDl0YVlUC8eVthB6p3HejxyQRJaj
1CBOfRQ9cWEG4xLgVnc7lbQ7q+hDo2JjJJb3j5AxnfdSvwJxneq22VgW5h8HcvyRRIfAPTWnUONX
V4AfyUS+cKqpnJvTrjunRAEjjS4fLtyalqJoHdaQySMFPW9un+s5YcF3ykhVwdgKrzrXmj+R3r4D
ASTE/7AyVNP3+6/44WDY7WP4jjQhAH/JZdB1+bGV1x8of957rNdrlg7fNQ3AtQbo6lttdaXTRDyV
F/trOgHRrD+tJ4n/ufoYQyJlmWpn9SG01p3Rb9NoVADnz234mpnN6E6Mu5IS2xaksK6EGNj8SDat
6WpDuMAChopXBmLqDn1ConKBvfyZgmczINB4TvDATpuP6CSHnmuWR6qK+qlqq0LqAm8HCVR77PoD
g6Z0ncXaFRNQY3KfDVVAeKWgNyyDwC8KdjtUykbjOTmtICRSLQzwsXQODtwttTA5CSwe1ouryZV8
AdvnTIZg0VvrX1YXHuHcEB+OSCvixq/gBZXYDEbXFQPbqj3Byg0Mhs0zQNX6QtqJHNOdJ90H3Yea
JhChqtP5ecVHJauJbM+MKjRRlDoUBupX6AN2H4H/DFhIcm7C2NnBJCuGpKUU+Enl+Zsl17U6HprX
hs1QifY7YqoK1QPkyrya0tuwpwAbcwzbC/L+IKaWiKbdf7qgoMiVfF7UgWPvZqtDcjoy5sJ178zY
2P03CCV5XYlMoua+b9M6t6GlmBM5z8qgpT0JG6zHGs7q0bcKI7qYUhYvikeZ5JIEke4FiCbi7H7n
Du3BYt+LYIkRlsspz3SeN4P1ICUld8ojL1HBqvs+w0G2o9tb7dNzhByXEzyVpgH0D4gkljWDMNDa
xdP5V2GA+rKbhVuelpQk9mLKj8JqexzwjxQEcbdw5CeTHPctUxUS6w1hiWiyS8XyCWKvC6GW8qiy
w756B08LuXC1WOxOhirmi2DyuYWD5V951hLFgNDgiIPMM3GK+8wNz4dDV3XSByQikg7qQANBja0+
cUXetoqKKl6RnVTy+aZPjQS6qD4VeCYnykl0mKPQAXS2mbyZ64oI6ShxJCs/Xk1yiaUFk469Gzcy
f2eHQ10e5ncLsFY50obxBddW6ZKUJyP9ok58OoyR1FTX3Fbb34rGZROtFYqaJNfcNw7fobDpGIGD
elwz3Qu/Lcxww/NgxuEPBs08Mx1O4D2Uf3nFWrw2lGh5RzoqQLGK7r2dY1dfCciaJUNhZdxH4t9h
YdiaGPgo6WD+J9XuDugfQO4j95UKdd159MvMddZnjP5NFRFVhJTwgGMnMFBA97GTXGFx2leocC0y
1RzSxZeTrFM+8afpnkH2NafnmWx6JZIFLvtqzAyB6jVYaEtcKADdeSn80rjcSswSK10LDEUL0mYv
qlFNu8oEXZDrCY9iisXAqwlOdN02kMUY5Mx0XChRIQI3PmCDKI9X3wSo1THPbPStFrF4aHVGlwWD
BiQJ56sGLcTnsi1bIIfQjswVIZ0gH2F5XcxnARhXL5Ov7USYfnW3YsQ+ICzNZj8o9ulX8r+7dh4I
uPZdpt/bGev8aU4MuEj4I35//dpf3kDLcgIuK5TtaeFrSGh0mXBPCoSJpN2MxesqmFWYJcUztoJm
kbFKoQpoG2I6e6Q4LHAS6PIfbMKi8ASA/oR+tyG29gvLh/XVCEMcGoCm9x9161KYUS8gI0ip6XxL
0PwNWrlQ63HAhzt/2iIeFSAGFytAASmLQrnnjpC6CZZN4lXhj++MXNWgezgU1qabkkn07YjuRIyS
DyVD+whLjMrOL+COByrDCjDSOaLHmXB6fBq2/PymDviVZXYY2LMLwwjgHtMATRywclwwJYKL3tKE
+TKbR0RELBHMX/EJ3On+2pvsr8mg5WTjIhyQ0Q4/cR4mJmRRKO/bVcNKdW6zKpOoHO00UAzPGLfR
mA0V7cBQBs8y5oDmJY8xcHedA5ON8cWKIoL1OuDyJocMifwfORCeyb3qbKcSB4PEZVqoi/xLWJue
RjWo/TWcEzV6oxX2+J347o/6wj5BXUuwpU2u5nIc65kVLyKdcM0+M6rg0VO7Pg9ZOu4+JEcHQyBW
lCxNvjxMpa89+PockUDrKH9k8aJmeANL3rsg/hVQbysDaokZXzR5fBAMMrMqc2LpSlmsF7tguGq2
FSRSxAQCYhcnibjeyLgzGOuebyKAiO0SCdqYgQZ4rSHo+wV0KuzqGxPTJhb/G5MvG5P5mfxwwUO1
RPGLpk9rfSlM2P+AZB/aenTiElaSlNI2pgEbgOvUF84MHRKMyu3zKDFRjLeZjE/7x2jfqpvyP0RA
K3RID3oRvb8fSu1EjBsIQmdPDwDQ1HkBf4MMs8s8Z3e69sJwyZI+aDjgNBIGk/hgUPpjRovsUjpr
5D+J9yGh89eOfFHs0obDpXuxeB9olkGFWrrcdmekaMTXEF3sElYPsKWqfJ5u4zjyTHhBAn218AMm
fXRSm9JlShbpl+A7sQU/8UGfxbFMb0v8ltDzmA8M9qtyn9pFBL6Stgs8fS8n02ScrfXCWkAsSBnj
+JN/IeioU+DfgtDMM9CaHQpzcpVRFRO2JRRJikVIpYo0W/UPFEMqep/w8+WzSdhTZP4eFztLLEaM
qQRgPDJtsWjH0Y6VwlE4nOyN336SVCgT++PqySZBaFYtn/0GXgaJLZEHQHLRSEbRwMzqMOATF/Lo
Hymd7TzZRAiVSLcGX60ZDvYreMekja4T/6GdesWhfgWTFf9pvwq+T+U+jvS6Gj7ObuF+2yTF3Qzn
bxthrOHW2Xa9gnSoIs5a2O8YKLc9vrNIYebB5HiyhnEC/QKoXI0PQvBBojn2kkaazxMb9Upuw7rM
4jMC7FgZe0heeF/QukZ2spr8WeIyumDVUHe96Q0v2wj6coVwOqyN4EpLdGwfvNr4rZknJ4ivowT7
A8SnuEloLnBR7xEu+0DRQVTTv5JXEeUTdfY6HxIZh/sUw+r/U/r0EEMc6ke0KcEVSqJSY3CQ5KeW
I/3q/cDTbdY89SEIY++6V2yPL03DhJkqSjDqo1KRkROJ1oCtd7s8huRe/1OYeuXyAiRMU4ZAY4Rh
s01hlH6hMV/IrVuS5nENqTgwsK/tXprChdTVR1AtEjNowhkEoQE9w0eHCh3AYQ50eAXyfQgaNo+G
U8bZwM19b4WGt6FSg25v8dTTwaVBl/0s5mqmWkp/lnAHtsleRDCyekP7IJdG7sDt+veP5HZCcwFv
SFrPJXKa6v4Mk9TNNHrAqehWn5xa54ObLH8zWkml2sNOa8rS8/BOk99AI0x2c/494xMeoBwjAiiN
8g3A98x1nOUz64qG22Uke0oeJo25f6QGxxrPf8mcDCBedjqzAdagTZOolY1SCUZNM2W/GNkum/FQ
ohiinGRR3IK/2V3BWNjlIRO+0Rl1QAUlREwT7J07yTzGtotAxZZXlaa+fBW/+4m3ZdDYo5m64oMx
Blcnx7WLI2R2okBXP1bKruuKfhpZDZ4WNaBQhIx+EVGKPrxIXu7gn1tmxi7wjs/RUgmgejT5nFt2
Tc0TJBTMBn4ae27FH7ZFrVCHvCrjwDr92WG0z1akA6/kvNhjJmtz7ezCB6+SaI3xHIvrgIVde87k
X3+yjOY87Av1itb+oTo8OSz5hVEAJmw2vsRNh3eLOdr5AkqDNSlBf5hDh0dl7ycD4H5snhDgKtM0
YuGQjCKa1MQZ6YTZa+ZVp0Oj6JS0l/03bqCVsW6H4CnseWtptn6Le6d1JK4eJZ9uOaAbC2ncesPJ
0mABDjaarMtqNYGfPVvd/Yx5eqeDYrWvRxkBYiv04Z7a7sDB8C33qYTIHMBJGP2Zoa1zI7TMOXxX
34fX8KwLmW031H0Q6UZ0U98yUtXD47DcPR+s95jOj5K0l9V6fhqMH3p9nPBeYple/CPoLVEIHF0l
cGXvZDEJ39TcO+YjcECmzsxMQvtzojo8lAjaulOa7cWcnKaKSHo6G8o6VE7N2vmjzvUUzCV1+gmx
Gn/64XDKeRU0PCn7E8vt0TztwZeybUUo3+m4oS9dF0NVRC3U52EvXYbYBnfcznj3IaG/SDk+d8/N
6/805yktYFqz0whZuIpqnNLagR689ehMYEJufo/CNhFTTE5j+lkiNU2oY/DQjkWKPlVLuC3lQ2O4
xCJqjOVMF4Ig7p8i86O5/EJDQ21F3d7LNE+1HSNMl4ud+jKFul9lSgY8zFKYowMqHFRqnedaMFRx
wIRE8Q87m8JFMTkC9pFT6pQlpdxBxm+GlEjWMwgg6oYBGw1Xa8hrMOUDZDtUir7SABeA2n4RKSUq
oJ88O4UcX/DpxzP74Kg5rcixQIsAfDVCzGf3PAFkLqMt5J3+1XOCAJw77I0iza2DdUroBT75EupY
kaXLJ93WR5m1njXL/IV2ZPcHSsAJVqRKyfTt1AV8SpNt5mbJGCpt3btdYieReqbzWEK3WrtSDXzZ
UT+jZnF9LmKtp0wQE8J7Gh1XbFc0DUJraB2Va4BJHJpqfbt8Lm+IWug3NvsUhKblHaT+XRe/Ah3g
+2U9OmIzr4MPBWJOaMDT4kwBVQdH3jD+ipxMvQdKk/0Wbjv1h5QJ+ZQeVGklC17SzQera3n1LD0B
PL4pmVJok7HNVHyXQMbtqfHggrzms+mJrLsyPZOZIB2E3sbpL5LvQlGs6aG2hMlGzdhwT/oPRwmo
Q3M5I4TQ4yyZzQzZ+MOlOFrTuMAEdV0ZC0M0OLj7HYp4nK9n1qimHyYHIr/A8jlk0df919DpWURc
2FWjt9QFjgHQ+Zrluywi+l0HJTPKuhyyWvrADqXOYyhJYPbg5WK6WSAns6GGVJPWSogG0dWFWWzD
zwSjnk2ZWa1QRKf6cgUZ2vv5UpZrmJ1PYhz6rB3TgFE563Usqi1d8nU9r9ZqgZWKUsEXtiz97RDI
BFwRjxkZtqkOU3pu4PX5bws8cWNaebZ5GxYfloeAlIfeywn6/MTNdG9srLDxNLT4xQaaIRMIiONq
Rj8Y10mctrt1etL+4H1rZn/jeWw3/CYtQGhvBH5ly7q0TDZGQZRLUoE/PX9xYC9nc8CscLXo2G5J
JqTOri9pJb6r4eVU6q0BYmdfjhHT573gm60ZyuriICGeqAEigVPvjQFHr0KhE9RIny/cjYrd79/d
E7SPFeQCHjeALolI7i61m6cSlaVo8OrhYIa55Vij6ec7dawjL30lAqNHxYILtq7GtZTl6qkzW8mR
++2LS7Uva+ejLjyiAUI8Lyh5PuVWZZEqJ0VPb8UILLAt0nzchQrf5rYeF+KKu02SzBHXP3dwXTEp
WJjBwhqsK+48AsLrx9knpSCtbX8N3kWvr2SMlpwIrqK/Dggj/dDqEAASoqONJHQwSc65xaino+vU
NHcanrmVPU5FF1PlLajNpXRMa+6wffPAlAsR8kHQ4x01vHv3ri3qHaKSD3ol/yYyhpgwCa4vWmIu
pseRwB3vT4RT3RWsho9VPbVUAUcxvrdVKoHGvfwaf15CF1xew65UWDLDOCTcZSt3TiXOTaG0IjIS
EhHf1K4VzInyxrkx7aeLCNrsOts5cMl36al2WciFJEK5JaTYpni7jSnDUCkA7ZxB+PRQMNQ7S2f0
PYOYWU3Nkik+nlpfpCV2/+ihc/EUBNxnz5UGXfXMXXk8hokEiwJmJab+sIGxnjePryLJRiEpFU8s
zGrInya1rcXXji36xBUipv57+3QlWPU4QwdE8uhmHHyCOVd0/M4LuBy8DRN9mPvnsRUsD1qiH445
qH/KnLlR0szVgoccfEyjp0B7lFRZOG+EUGK+5XGCcw2V7lMqTf2+qjApjbc+ZvvGnxmSWEPp29Jz
Zp3iTrLaxL9hHpzApsUzRKkWYk+QaliY3ZrhTEHXMHtD/wE2zGmh+lduZQ/ZCZ6gY+8opQq+l6xk
3mvxxme6y8n/o4UFbOnff9MF0/LRkCnmMO25OS3PGA+hAlKXimqMEpo4hgkyyAfbHep2El5fL5zd
Mkf8e1MVOOvxEzkpN/LQJbhA3FTSdEe9AlBhw1vg1tznAVMHz4jWCk15GrKH5CCX5c4W20b1h5zE
Gfxxj+kY6uA4a88tCI99F1o64mQElHRUkmAhiXNqShEW9l9pKxwWogwGuS/HrN4YsvVTS780bmDj
B6lrhC3sM5QB4xMBZxhiSsAW2mDRCoaBR2IvNh32dM3apHKzWsKf9l3YxpM8LpHwKYysXrzIHQua
uj32ziRuua3mnj0lXkCPQcGSwRoB3cAVk5w0a0qnPVncujTvs++KOG3AXpvTPRz2mWx/zYau5e+/
siWWgHNihwhuuWGgJ13EbWjBZvtJrAQPxM8VOYgyMCTP/guDUoMCYjFLRaJLD64+6nL+z3uT+ZHx
H933X5gFeOHwNVPyypX/98jV3YoXha5MlVNvtkJ5LXr4MX4xQHl9lXd9NQbo3xa1cUb7A7MTJnzi
NcMGaosLg8OnGCNDjanqABxpC81I1ISlfWVXOs52qsW9y14SW9axoypvO3WmzzMc6M9yEYBbg/9T
BJplSya5dzvRitoDHggrcBqfGQDNJ9xB6Q4OmTWqGdk5/N5jT7RtmkwaiDhayTBjODFM4LOqA9gc
BNmtr9hFdUSe8EBwzsAGWsY4H8bFpD+LOFDz5/SaSAMSM+EKfcOffVoLKBBJOkEfi7TN7WKvk3om
cBWopgp7Rkmh5DeU1zuT2cZ6RLjk/MW1d8lIrUdHQtdMwfmxdGXICswZR045ur/TA6dVKWUCZDzq
hl9UmkpLmjky7ALMRq3IcGUAMokse5qMCpL4sxup+LHEj/66uj1cyXL3mG4/8pEQFzKeQGxUUoAd
P8aKd+rnPLOJ4C6ifz/usQAtA0BFLaLNzvlmelvIMvBadkLwOWlgG4KZGAVKNEEtE73CDN8rdVce
tzZh75tRbnX3p6C+rccaMPjOl14mN1B/wMEmjLbIrXKxqmfhbl1Fi0rmqIdif71e56yKEIwlhvaK
8rUYfJAnTc81t/Vrzu+D3DpeV2IOVTJsfsQ9XjrMeoUddWy72nFG2HOeC5j7NQAtPKA1qEg+v3gD
d5xtoZ2vFMirPZypezEE/XbsJGdmNsS5CKWOzQhN7J9Gh+1o63Gb7fIDTnjp5V18UghfDVgM2aaj
be8rP87gOygDMqbDPc2xpTqqRluY22BKFx7dExHCnjFAdFeuwzzCu+W20u6NAOn1LUpC0wNnmjss
QQrS724OorBzAUy15djKJUzFvQzFc9I4WP/okoa8ZblQm6MKNeK62lFiO1WeynArJDgtD/54eD/E
JRF2e1cQHP5JrofxAl0I03XrN7qual5NDm9NBjpUTVI+LVbFUvj4yA/0yAFj++RtjZycWQxoHu9z
GPs/D37JKTE4C6sFKiPAajCD8cuqqHWJabRMUmF3Gb9xgY7qn5D9xF6LYSNG4BBOpXpxmXrL5YFc
HFLUcTULlh3XaV/yYoIL8b8I3dw1AgIdHdodOMp542eEt6whfy+TnPsytnPYTiAJn51dr+2rjSCh
p/64RRuAP0NCZTDiwgKcsoua5eM0KXrqEtCyRceACubzBLthrRVJpbrh50VmvbZU+SvOuIo7lZdB
BefZFrl5h7nSKBJQCduHvVgZpKD9V98yLysN+mwrc/fjvcRiXXFPh15KzQkfdZ4Ckj8A2enzJin0
h/VKZv+tovdittd1jVtGSrNid7pq20+BWQgTm88oUpkPtI1R6nk0saFDOlWm0+5HrplqdV0xAFF7
rDaJxaomiNWgFp+86OxzVJzCogXq48+tYV7Hs+fxg98xIVhESvwcyQQN3xXP4N+CHu1qMiepq9TA
QEcomiD03MKNnB4d+wXLiAzyIEu6m9MdCwwYv6hLFPm7Ws1ZY2WE8MiOtxkam8QD5ENwUlHmPqbo
7bPTc5PxaQDvr1UPTi2pEP5RYupDHXX7uwoHzLcAint0mj7476tN6yKhNg0HYZMVdEi8RqEs3pF5
9rL4t8p1Efh7YLehWHRmrV1uGYWiE9rX1/5UnfcyDf1roCOvKBw4+IHRTmwwnExmNp0I9CLkpvCn
szUaIYotMFYeCGzXGuqZmclnt1cbsDt/IRaDAAIbogSKfjfcZao8uQKSogs9j2uNCafqSgG6irA2
Ygz/xGnN3AKmydxOs4RTjE4+mLvFZccyqQBHLCeq1S7Nbk+fXZwQF5ISbjHZnDokGE7T0uZfO2fF
J/m2jk+5AKJ0hrahVwv75Q7VA8n135kGsoeBTdOG5GkHq82xEh4AyIRIqs9bnSCWGJkvDCR7t6Vx
L1TqRENoLfvzf+CSbTW8ZnZUqCxjiiCV94lY520es467gV0Q5myxm/UnExQinUc+X9rIBaOz6j2e
OJvCAtoepXn9do/nZSkbEanR3nnK9Vx0CiRprNKgli5sCyaZHC/G73E99cZkkeDGpgeCPsp9IIHB
/3/Rxlzyay+GgQY1zlLVNCfTlWKct/zkO716z3Lh2HeYLSBqaMkA4oOg/hCYEigQQnr8aUaz77iW
PriLAW0vVSgWlcm3xdwaFvukkNWbigA9BbjXT8l3IMC9CS8BwSKT7foAMY9i2ipQoaYPGH8ZrnEA
B7M49379r2knkJGVVRlohu2Oc2am5fsDWwNxx1fU4xCFlTiQhyl2iwQ1KtBMUOvcH3jAsyJPXVn0
1uCHWL2PvOwpN31OpCn5HMNykMCrvd0BzHzVcvImcPdAduHQaX7UTHN7fp+oKb2WTQDbnO5K7DZA
Itkw/gmTyMeDTB99Lo0IP/y0P90ybW/hqypVWb0y33arFqc2ULEOWJS49OmqCuvtHy9o6mn4WxLf
ek3JrP2Ze61o1tSvOfgZ12PCCycLGXJFSdZACmpBLdtrYHrgoEP2UTgRtW8DufPulLt/ZVyXy1Qg
Fx8reht0leqTy9OylHzwByB7R2i7TU2bniu1YjmLJdN/FFWlNEX93drsLHKUQ0EOBF5A8+Ya9eHv
QWbfKP64l14xLZx4zxc/n1/eKaDXXc5/Cho+GoutJM/faNf8aGeFnkYFKyl0mzwh/C/MDi3Fe8fI
yreJh2KWjDL+E++Ow88GJy07wCNoSrMUNcGPM/1DUyYy6GrNnZ8M9bhSve7VXt6H932SrCQUVOn3
9fM8vyZQHU8z+xWgE7tJYiz8DnESoljM5yG3t6SN+Xwmqese8IDgIvpX3MzkhDbiTj0+pVywhK/L
E2RTN3gsUlC5nlLyzgT6LUza8AwFq3OY2uCWd+wXywdl9rx8Ew39TlOlOWhWi3JQysyv+ZiQzzo+
W6ZNwNCMLbkuM9zIm0oRZWOyrZFtJ8ZMCGhFx1HjKgykjiXcUiyu5QuqOhMzd2tOHle0P4/krAVb
GDFhMZ613ODRX5bn7GfMso06NuxTbR/kgPhWzFWUwTSEaNixFUaXQ9N2S48YhIvqJ6Cx0YyssCpo
LYOhs9T6yvPMwCtr0yujaTeanCxkuyiOfbTltDkvhztuP6PZyo3kNkt2pJ4q0JSMiCAycJFSNbEX
KMpxy/aTm3iheBKbm/7OJb+Wi6xYbZt51214aox+grUJ2iaP3CH5hE4xvggSGREqHwpIxgBMRccK
1rMXqGA5UThfjkjsiTl16MKHeZuFKfp+BNph69wn3s9zG5fdpx9bSx/a2u/fkb8OVAASfEaJ30Bp
Jkpggof9fLX3IqYP2sR6PJ6rDbUiUm25rn7UMiv3mubw6zkPZQXrD41m4Mw5Ct5M5R+ypkRE2MKM
m8U98kI1zMbfxuWJiicKfI/fE/Y2Stb3uSR1Kdws5TaQk5dNvcNQxXaHGVQgHKjMCOa5GB92HJc8
QETB0VU29fxHcQ8CKZyhXtj6VHHjGrNgUDPSq7LQZl0unnegBs629pDZMuocNTcMiVK0SQsMjz2v
dOGvv+R5XYJ08FqdGw46fwconcsOcC+Z0xAFHk3OUjoGdmbrFdxcPcjB+2hEXepjn852ekJoBZcp
LPvQtUWE15j3wLBlF5s8cG9xsUFlodRk/qHzaQPih1Yo7O5DawwOKmghMBELLMF4Tm6ITx2X6ojP
AGMGeSQBUroHLxDZUuYpAkorQUaURsADN8scOisA81ashD0FW2ZxgjYje+p7luX1KXDvB/ohtycg
THw4TIJTqValUS60NNi5ugkMRQ/l+C75sKfGMNWLMLgPblexhITonNz4U9Gfvg6KSL/kMlPO37lu
qCvqgpz8wemRGQGwJSDDsrSfA5rTe7i6IqcRCh3J4WYYhQx8Rl1curXsBN5K1SJPgzGPcRWRCR8B
OUI7QfR8hNes7beMt0cm/Kr2bfWSDwLgi5DVtN4ZUZldj4bUU2rO8HDvHzT8Wxtfi5p9mTvKuUwD
m+mFjr5SYJVySrC9iNRO8mQwpwcZidOL3P1jJpzGhON7RwJ+7kYcODwOt17MandIgYOfawzYWaxc
a1gW7R46E8lN2MaQ2+Dkzd7h5DaM6TDwsHZcyd6iqm8GgiJbGs2fSzfmIHWvXGZsC73kq0MeYz/N
8FKB51uHZC0RCmi++sAVJ7y8i4DCglLhlyjhfCoDQ37f8qeCz4G1SWeNXXynaPbyyeKvxbz0zKhS
BQ5L5DwYX43AAgKbDC74Xm71BwIw4IULdQj6CfYdsP0Editm1hzMR1QJ558Ck7eF6VeejFEwn9IJ
cVFLBoHyP0da3Ydu2/pbfEVENmS1l+rFXL8v4q/x6quWHY5iwAEpO8VSrPxyJrGC8hPwONJYPfgR
QooUXjQZBSEb9gXEVN51huhnxHJN3LWtAgNEvy3w22hZCtS3YQZMMjolP3RnnxBUo/0wNqvEeM+R
GV1ur84MHisauH6Nalr7FWXiLBqAZVxGOHW2vs7KXLg08P21U0I2s8Qdp3EqYQ6EtTFcSpoagwJJ
yYMn6yRadWEW2HvFOJv09ZU+dJk1eM9Ba9TxtAbrm+m3R1Kfw29B3/dFpqhRBhJ0DbXoWKqyNIaf
jUmlYFVO0LrcAQ+X44ETi9bDpAgiss8kjQSJ5SIbn8egXSpHz3AD/F580semkkl2RQST8+CQtOMl
JK/N2pF2TS5hvZMM4W9K+hvps4VqB/sdy/Kto7TGcvSbB1mNGWZQJP4P55vkWr18QjNd/+awC1QS
/dPsN8EZNGwjyY8nplRORgd8zeTvyc458kR2cXlSmvmC6zVMDufBKu5vPVfCFkoEk781XN+QkXbH
POg1cfGAKLM6fv3C7/ShcPoHdFlAWBddkBe7gn23QYkjadWCB/pTKKjPetGsk1/QNJYzNWx5lH26
zXr59StUX/9c11hrA6eCOcIuWwZcAovGFVz28ZdZNIHg6kmF75F//DYhkAbDrwFKbl5OUvxokeTR
4lksDR/B37legjTdXtuxXQfyr8CbPZXdFawBsgQhCWoEhBYurzjLbOXBugWQoL3dpAyNhM6HIr9L
HhOJZiND5tjur9BNT01Yv7RZJt/8QUDeXj1Zbxf2X/Yzcbbk0yFNzm9+9FuN4HzPBcFOeeR1fT9I
8GNO1IWiQndAK14fYpl1NJrKnwgOpaJYJ0N8c53unqdlHTsYfVF01mSjUX/KblBFIF0r9uAn3HTq
4x2QHM2OVU8CgSkjbUr+boYLztpr0coi8PzMXZQBPjfWnCKAowGzSMCdMz9D9TOzZRuGSnydbkF+
wkgQKjCyrgm4mkIcrfaIUG9x6LYyTtHTJj64aNVd9LA4jpurZH5E/0HPv9rler5U+d5zsPBMJ+Ro
q61K940yV5JKk+zvnxqAwAcpCruOyq6Ip8UWWIktuFVmMZd0h1BI6PzhqAxZgL7YWjMd/by/KlAD
fEZWH8tVnPwcL7E0vCEOorL3QdHjuSuq4RRpiPVBYsnY7/sbJG3YWkZsRWeozaxESro8eAgsgHZ9
13Im4A0/R8OvZil3TLdtxydfeXTJe5gouvvsxaRMPl/lI/w5NGiN2FVN/cErs2nIoannZbwup1PO
VBdDitcqjvaeKqBtVHrFmWNaOkfF4cL04sAxjXOwMe1eJdyoLfz6dJSof6ye1cXxh3Y0M00Gp8ih
QvB2+wbAeQs5P60+VGn6k1lJz1KgFgFUld2Vj8lcaC0uahYn11+kZA10g7wm6JpjSk/3CUnQUXwC
mMFHDE7ZZnPCVL8ZOOOp8nnNSPhal310RfQHq7K2sB8CeJZ/Mry/CH/TJcaxpShmZdWCqQzEQmGW
bgQm4ds5KpkDQKKc37fN/Dx3M8QCaaCE+j6AIOmEsnaSLx2G7JL9tasNbgFSNNwtqAUPlhPbGJws
R5nP4FGdr09nmtrO/4SUnTjeit/vWKvngq/3EAEca0Hw4pjKVX6sedzMvh1IanJejJTLzHc7iZP2
MR3y9HHV/8ohwKuTWjbPs7y7ueIvt+TOifnhWkbDGgKl+t8Kh7rKv4lJOMLylHmesRE2LzaW5cnL
I/T9R6mfb8tMtGzAShXPBmJ/3sfZ9lrmfkqty8gzHGS83BKx2Ea79FPqCMEDLCWLu9pOxh7Dc2tT
Gp9MYFI07AZwl6uwyfdrpR5UL2J3sEOIsk8Q+loXPMl3Ra9TQZVZYIMdRqkBNVjxq5EHwutPKHHI
a3erAGbOZ8Z8MfZ6IxEbKhWHTzgvDK4ugTU0I/kZPnxItD6e2wk4thX0Iu4GDhQQs4ikRzHFTouh
8eZPN2nd7pUz+bftvj34u/GmqkWfemA9c5h7IVnZ21G+Giagcn/vDkHpUgdABpMxu7sPkTJQeZkR
MYxCdFVTrz9YoxstfmqRBHl3nROvZho4tdbTZWm1fsBPBGm8JABiz5G+BFn1p5aCa/wZq8333PPm
QQd2zLwXnIAj2seUW3eNGEV+H0B3yd+gAJEisJVtneZZ3L63/G5NjVi4R4/IsgK2IQviqE4vfULS
F3d9j5ZriJTZQuNiu9P1daguC85bqBPySDmqN22b2X3nAfIBxp45nl+G+vYlCWgJgceY7eUgBAh9
5L3MscIaxxSYTxjlqzfmVhwluUXjKvqNhItLT9mr1SHH26DyWUv8JIydCh7CXJas/aex7dgnGuWQ
5nhuLV4XJfs9O69Ee+hLVZm0HwUQ4BXXOBUCNMb1QiQPKVrqr5dZnXtjCf4JsC641rSlQXh6owmR
csI+LQHnVbeNtI8yBF7kMChrvEb8ZrT65IDzmpA6xzgaU749TZKr7IGRO69f5VHgvYRyFnlvS7g/
jE7/V8vVo8ARUjzyVKpJ/yFYULyc0TQ+ccJ34jdz2PBf2pWWJSVHKqmJc0zisQHYk36IMqk53iPo
8WCqNbzmWP0xVwhUIlqT5BwtUqlTePodZ7TWO0VMPlJz4d6fyx5Xo0IelAH7mn6zSLqbYVa9NpJD
CmX3F2O2lyPZkhaQDC2v4rmMGTgqyZ7A1sTmE8b9SYHR+tJU283c7KTGenfv3W3Yc/vmXwXva4c5
dem6Hwha8o+kttJ182BeykiOFtH5xCDJKgFmrRnYC4Wdw5C+CDkGANXDjrIeVXhEgQYzZCGeNGGf
53pPGYcAp2++Rbmw3PsM9e8vUaOgB7VBLtVwBSztXm97KIjB8YNl88qdAx9/IpCDGfzpKWO2l1dV
fJM6exWAJA8VnPWz27ThZ3OQ2Q5Se5fDR0AmQjMB0WMBjmh8qTBCpUcjy/Zl2oY4nwbKK/eBrmJr
kgvRdhE3WWFjcMTtbmFEuRWOXs+kmylSv0CtV6Y3ATSStnVpE7Ya/BJ2KREQ+sZ37aZuhHHo+INl
srAGurBRMt0hYG9IAozqHttCLQehKPVWJXd50NoY1wLoX0Ei9skmnqKr4dm3tEq9qMZyK73EqFh+
pZ63UXWR9ctrFMy288dVFmthok+j8J2+9Eo6Jb3eeb3x036zv9/5o+YP1svjH20zGbgVW65Xdxod
di5H24fgen66kArvhTaTmq3U13ia0Asa3MHUN7OGwX/yDiFSo3zWxox6xRhPz3uE8G1MI9NEAShx
GvOGUKVYYSar3qemV1fOKRuzurEsMZMLqxP4SLx8OrQCAChM6+uf+Aos0gDWnpw4AQkWrmWhC+a6
cx6VyMFvECVsGMUHOlNZr6dagk9MCwsFs5PIOXquXNlbtDT+XyASzLh/ghhCgPjdBpvXjr/HY+Ke
uvljjhwFhB3YQFO3Da/bqUn14pAELS1GVpgUbpLAu3N1NWo5pO5VD7r6fdhKc9vZjQYR2szQ1j28
6JBr8viaMx6l35qMMauEeBLT3UWqsaQm7bLWc1dFY/SJ3DVD70cFyo5hAhtF3wO6VZrAqHLaQkWZ
+Ya5JMhiY0pYt+11xR5dXtDlc9x13OPdtMoedZhkDrrftQsrkPZVZj3rs+L4vynn1uNmHrmNTONR
TNPwA+wNk5q2ckNelGrZl55lAFv2BzrhLGpXdnwrxPgHdl/89tPCKlmghS3Cm1yfVgWWA4C+ZyIf
3F3hnKru7TExp8hJqziqyaqI9ZR2QpflW/Yku6grgnjYx3oUp1S5FuDlgsVLCjDgZ1dJ8f1p7Nny
6xhvefDWAsTJlfnXWJrt+DauL2/gZUZP/Xh8QDsLHDDnsZl9/8FAplt4F6W0tdjvI9wrp32lenVg
hGvkrazx/T2ISPotEhoNCqTeaZ2hCWgWdJxBLXhNp0esAE7c7iKkMcBAuSLDbJiK0vYnCuXU1H96
/IBmwTNCS3b+p3ncYkpPc9P9mFOjv8ly+OJvnV5sraQtjySNEbittMT880Z98PdzHrEJFsZ8HH/M
6pAn2ibb6qLWLfSpAqdzwqo2AmP0v7wPOnNZA6gpKwx8AExnk3yG9C6tRYTWpddOZxcg0tRzTdX7
lkuQabzebaKIamrv1X1whDY/ubid6P/ug5tKV2rcgl46UxdTBdQOMSpva0FGXbF5n5Mp7n25wvnY
frBN/tOS3Heb5KSzZPPDSMk97U2wnIKK09iiVUX+oICDKChje7OG3R9YcKJZLpfS+lRefzRhkf4f
YEJVT036Rb4m7/LLXzvT6Cl9aOfbCHPlagPzOJmy5Enc2cP8EgO8k73VwT/D9sruaEo188l6FdUc
m+UmADjwf8h4QPyvRAPeAtEKMoiFVVZn06Kk7UTr/6whZ+o1f2KcIocW9AsnetzCoPcVWRVQacuW
NyZt87R8/90sXatbKIx+gAKJJPQuUcEV33B8qyX30hSFr2llDBsNneSUBvqaQ88/gV33YUxCr33W
6mF1r/TY2Z/doAVcrJcUPy/CYNif0HWfZThV7b+mtRbzSQyKAk+nCiT2okVFr4B4U0n9Hqos7xyE
AiTeHyDxPq/DV57sF6ZYFCA8QKfGPZI7EKu4UFJclTpAcBxkNk9qsOJrK+nBvtUQc4cRkaDR/k5q
mYtWNd1GrKSBSikSpdyqj5xvTgijcRwXkbwD7cS075qBccCFMatJNk2S1frt0krLjZPcNgbO6Qvd
1XLLViAkzjc89vSwzprUw0XoET6BbLf2zbIavxfNg0dxjjIY14zNygbT41jQlRtw9mtNNgbUjGIr
jUsjmtxAuXTomjQbDMhmNewpGERQgiDiLWPsw7KaLXSiT1aOcNfAl1uV6N9ZbadCBIceU1HCLHM9
nq+qRBVRrOeJjsrLI4Y1HFQwaNbqRDUPElYnHHRAxCW+9/DNq2DGvOuOfgQSYwBfc+Cy/jv5dItj
geDlhKU1qarxKQzcIAEHLrxHGYMRmNAVxWGsBG4Nb9VyKAZFZweYaStlOWJXrb4mWMM9Mrffow+r
szghUrYZhPsAe5Z7cGLcuYAbanbZ9BGRCrXyac5f261HT0wt1fYhXH8qmRmqScJyZU8daArYPP0h
yjYB2pFaj2mTKba/ab+8UdIDNjCJNOrc4Kx3YMkE94vG4a1sSsz1Ichd+n+yNKNBu+U18tLfenVI
ziwlslyEkLDkD5w4iYtY8wGo2syB5JtWxRI9kD/9K4DdTQELbIQrumUDwAFvsiOKmOflm+7E+NI0
p58Ciz7n3jWVbC8cPdwldx+5rUTDWmZINjEzuNpOYoWnRWwtxoQvA70q53D/bvkwVBa4m7Xw7v73
05g0fSsKLfreSJKBKoGll41Ox/5DVSAKWOcULw+jRoSjjkDa5R2DycW/a53oI+soNYwnyhIQaPCU
aEpTTpgC4b5Fe1ZE/UzaQWEWtLHGEWLGFQvEO8kIAshd5RFchNPNr2Vn8qdtbZvQMe/86afGqNae
NBU4zf3JE50bBhK3So+vwh2e7HiQAaEf5k57X6lqHYSlVuO9FgWF1yjP3mHkHsUGF5ewLzJLQiIC
5pGmeItk8NPVwU+x6Qp9NIu7+VvnUKXjvQxXFzkCU/DVrC3+9Bz40JALxZy6oC5TW4C2ddcXVGO8
t5GVTg+OJfZ3vjGNYeeTvn55dwOMrGLzjkhIFT2n3GelRbkHLW5vHP+w0Nam6WfMb/AGhWwrcqHt
/wmMP+QkKTfKKf34fA5m3kK4IZuDRJGMXY4A6RBTEWyF/QFj6Unj2MyPMVqt9Rs8ikuHkHz7Z+CE
Xy//qUSF5xHEDVG+c+7k9C2Kb7F8A0jXYnBuThWLOv3F2OEFJHoqljvu12JBkO8k/Nlzj7eDXPZ0
0RmXMZJj+6XMNHRjxDU63mSPE3yNW3LCZK0fm+ERL5mQnUoic/ixdGfw9nL3NIngLXkUGb2i8CC3
1AJlFNqPH3OGW8xvjM9a6DLJa8nFD8yWRvi89fT7I4/QMFcDovOZCrh8hXrPGHU2GtaUe2TIJ0aT
66RzR++b1TH/pSpJfTn6bpymGNIPTrT9827KdspXil42s89haJESfwpPFELM7JdTIFIGAGbyR78G
v/OvCFWkpT27kj1L9GKNpee7u11FJ0h0Kv8H39BHZ6l2dEiGWi0/Ey6MF47cmNE5VIjqbkY0HJ1e
3am0dKil2mO9/22hHNJlKstl5I3o01e82ZU27XhzB0j3PRZq4NebH3wkCD5RzEPD1ZqyfiKs7Tz5
1Pei6FlrbFeofanfkJntJfvmlXh/RX36zQsl8KIu6mIzVhBZdshqw2CTilXH4yahiHbKheQqoyiw
EJ/LKJYiIKep6owjuM1G/HbCqWPuEuuVgOUAtVR2sV/hgFIpYtBRIAaCo/P4pNI0FqjyTEwmRKV4
vNG34wnTsPgQC7OH71VkdAtDiU6u4QN0/jflEf86s9V9EP6iqA9XwjJBvFPOAbKsxBTaWiT0ZhL/
nvmILICR9kB+zd5+vGsZvXQ9N+G1w9h6i9tk/g7fVP3uMTJTLvBvhiD4xqsM+TR02Is9RmFBzygm
zrwcRBNKGDotWLQ0Rbp9j5GNDXG6VW2t0iRI76uJOLSICI+K+4x+CTHcjFj/DXfniXOPWz6Qk0Km
gJFLO5sCqHLEgxYa+D6fb0Rgi6vArTAsLUW+0JCkqWJ1fhNbkA1lpgRi4+4lI7/nPlADk8jyiXHS
2MYvFSoIUjYi+cx419EuXumIJKUf0I9QVXzqgCuPcmYrYJ1cWUjM678WN+LAVPUXDNaceGkvWwXp
ZUAt85iLg093Tw+jgKx92RSsN+T9JEcZwMOuIXZrhxmiw0YkPRzK6DmOclx8sRy5qEQ=
`protect end_protected
