`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KAioFAHYTWsGd4iPoN3EYLCq7rWMGrnAFLwf700frKkumU6V04g7tUnOUEMvhloUZ2qovYH7czU4
GDyIleec5A==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a0mt1Ppgkpm3fN/cpbXYVx4/PJYIeSjmorcEAyXR5gEtq993YputQ/ou2QqdMuJE+itmMagqGTdM
i0qK8aArcH/TNv36yK7o4pDl5ctqFse8yUBq6hPp5U4DmuYJUcyuN2mxi9lMz3hNiWM5Y1lfDXNf
SUCkAWXrtYtyffZTL+g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V972bWpVqkmsPw3zJtGjwOKsiigUECZ2LjAMvdqi0f8QvaVvzlxx0/VjMWMuPEEj6LvgENW09mNu
46dJAjkFCUCj+nvWlV+SISxs03pO6rQNYb/m7ciS0t4mr6kGyfSU2YztpfpLqVrWbPpyElhoYq+d
HxDiTr7wMNRAOLS8EU0UuwIheKm8+6qhdJwgunf0fNS7+c9L87acEMdLrKEfSDB/vYfBGIvY62Fd
rnXAyM4suqr+d8jk0rIHnQ76oKFw2dGrHcHNTlIgFnoi2WBSBEL2C0yiGh08fb7s/FAEGN/zQFMg
7F+XmrAxxVr03ljZH8QuSI7CMhwcEDBiEqnRyA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OOn2aNhZ+qGR/ZfxbSNtb24omKdnlzB+Q8NX//Xp7h5+VGadmbxPLB2AZgZt4Dnr7wsCVg3p8T5G
SDXLBEB8rpWaIHEo2tICEA97mXHDcC3SlTyl6cDFh/A0jtb4COoXJ47KirsgJ8J+AC5oZ8eBYCKz
bUjbZ0OzmkQtV4bgqXc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
icNsF65C1PtdWcdDHtQj2ZUIYdxvmQggqKj5rSKy6omPkTd190o+czQZhd72Ldt2uLqFZ15k4YX7
k6qs06/tzEt+KPCZgr0/J7CHDSkIdVq0vB9ChpAIqt1n0MpsA4rBGabcupwQHga338nxLPFJ8763
SqmNY81A2y/dMgIXe3fP3E6ozmn07zDMCPsRtcEV4VIhUQq4TW55V8wJdC7pFM8pPTxBSyAhGUio
JWbYPZuoqr6bDv/h5Ganan2FkO+dnqmTmQZzh2Dv5kJIfuXuWb0PNRMC4scwSqw8dgOBlmkoKwr/
1dO8tSHKXM0JZ51I9tgENGUee7x0y38r8SzuQg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22112)
`protect data_block
wGv/is/1wTGkfr7+VrjPEx7wCvCe90eFxr4S4XTp4DvQm1cBy8a2OGvSk1dCJ/+K5jp3Y5SUsrDz
/3xbFR1sWQXRBhudMCxZgfA5kLnmXcUDF2ulsCEOnxWRv2+1vaSWnTiVhAQaMg7ScT3Kc/B6zQl2
U5NNk7zvrkBadrTnvD5sFgWQUDUxSuJMhKk1+kz7WiTmt1ZSaDbkGtEH7joHM2gWBBITqI4wCeUg
6moU9g1nGdJhpupWM9qweRneDwU6iVRDAL84emMHX53D3bfDWJkyfn0MG+o/3GcaotmEjx42ZsIQ
sD2paDWq9OOqS+GVXs1jWuFSFQztvpwu8oKBTThpvERvQzO8zgXnVC7cqS8D8kjZEBEVHn/KTZuJ
ySV90WobvM+YOXHlqTax2nXHrg4fSmGPOUnCMAtEK4eqEhyd590WZiN7TahuzywcOelzZTw26GAU
GnPYbTsiy4rHC00LIYWIMDBdqdOFQrCcxV37EM7F7HrdfIzsjfFMu37P6JJzeGc/xEwAKQgdG0KG
6Ejc6LXQfq97ddG7+UnUHcR7K6d73EYwuZfCFgn8mZtcgf5seiQdCjn2SZFTe6N4+Eq6CvjM1Dr2
I74ufZq5VcjbSyNd8APIlKMSzaLPtQExly/JZOWX9uP0Rz2ZdZeRGBgA6g3nB6CvNF30/v33szZj
k6xSVEEXTMpo7LC6TB+hmc3F5A8s5EC1QUTBQf+M18zLZofFtx1BCUAbRAVSWGaj5yF41nt9AnAZ
aJwHl0wHz/6Taj+J2JSNGRWV18Jad+Gmc6U2lXRTNbC+ZiNTd6XNYY2E2PUr64WlfM4twvKAe4Oi
63RpkJejwtjcMSaPSa91XuDN5ObAYRgIKKvYxRHEIfe+oRB3Yo0B5qHvZP00U5escWv4+z+sJmwP
SByYqihjlSYctFedoObIBTD2NzK3x/J8bbkZWqwATtWWF/gfkkBqK1F3d31IzD5x77YyPgkoEvbj
Yq1V7CPb+0kfzFJuuEZRy+S5n3dgGYw8JfWh6RhXePO+VUcCywKl+5EU+/MuLi5nuvE3R+kpkoy2
JXUNyqrwTVTznDqTbYycilOZSA4F/gKJNPJvfxMeil8KshTUhLDowQGjdaBLtV5uRFHOhu3PanV2
ymJt7o51e+eN056uU55+AQKutDVz4OYvqB2PFsUf2Wo9BpMeQ0LMHTV2zXgF/SnlX9JWtHrSAYXe
WIl32vUahdaWJgqOXqofsBMKeIc1bsy2yN0PA7Ftx1XpFNxb4dlNEOou5GkBCtsDge88p82+sg7s
CKk3crANzd96hGPHbNcIKbbxvmN9klBrCkkpG6eogEaf1OpLllY6J2y8u3u6+X5AkzbBVZq5bAFD
QmSBDiEeDFAa95s9i4xqQEzPWZpZ/wNZUcj6k1oo9jWfYuuTNyrzfeK5b9OcquQPUmLVrsrOIxEL
OD+TysflZmVVOlfgjg3TJSs8zndJEQPviKL7vaH/gYseqHacDf5mAg1LtvTekvXcoRKnTY/HZubi
gz/zUN9TFKoxJRIo3dyHqHDj+HYKzJtBaQDA5Zc19a1+PW6SiT21qelxaauvef931kpPG6V4A2rq
SQVtwnM1kcC25aLDNbi5q9I+YjhPLz3E43ImjZLXn6fYM5Yr4+nKSY5k8HNANNjBDbXgjG6Tn52k
GmASma1G19kIigkf/mQ1hmbEJg8O35ZN26ATWVVePX7ls0LgY269keQ57txgbl02Oee91riLKJeU
NTB5t1lwv2eTs5flYC/CloVJiyIB2Gzrm+tcgrfePCVMsRRYYUSJfFOg0U7rEvMKLsg3c2cJY2Bc
c800sJyryHdoxH5rLI2dOXeQ6uY371DImqrb/gcb1xIf82vQrGx1FZ6mgUTrz2GsEmC/V4GvRUKE
UiXQCCGzuD0W3EUOF1THu+Yctq/ieeTpjFxvSi4BFlawzjv10TDS2ycZhbYm29F2lvcVtwkxIlnC
2pYaGhqFrOcmKRNxZ8inSnty3cJZkSL4Y9YOXcsVX8bFNFFCOsDKJ0xngUQ2H7MbeZSPgRnQE8cs
Q/bfHEYWmWfrH8BrVNByuB9X/LIFvPqvlY5c4sfZNU71/fbJMJOJkx+q0NNtZD5Wci9CuJd/Midd
sI7MH1stpWA/ER06KCSq8cavLHB28mglZfD5cpdxsY194NeCv9VHp3Zq4fqQ7h8gCADI31gKeOLJ
7cAFlEz7Eqc+6OE/JeZYTTLSnwTPTGonzI/U4/aH8ZMZTV+78JAikdW42k3FWXX3jB2JpHAL63DG
pN9ltld9pookXJY1VlDCJONrRjFBU8xCJxPB3r+MMJmidiXuym+CiDX4zDTurTTN2AFHgOS85wGt
DSzfcVUmuEPijIkx+iCozYL//rVc1guV3bxnKRxW7CEElGt8vh3GpvuDelF5DtROBzaFyv1M9xWD
e9/6w6A24j93QrvyQRQQvCfON/Xe+JaqTkrmIbZaYMjyXNmEKRuT2P8AY+9IOqzA4lODttvkbkyo
OZEGGGZkLkaFtGQHjU6m8TQ1F5r2T6MI6+vTcrPTbKr5VrYZeaED16CcsyiXjxyloHPoqjqXNpeR
DqGki2r30iKJ9bBJv1IRbS04/L8H6awLAPLCy4RTyyeWVKlLt2TgyDwntA40MXvSZhaXra4qAX7S
r+z3udHajlcEFTpQRTH7gKJQi9oaABwhvageYbjaPHHlApysyzUiTBaLVUQg1DOj1M6r+8H13q4+
hnOKXdx6EdLr8gneUhT+rl2uXswAOvFl1uHZzrH0gFq3fjARlqXnsG8g+yyXs/0iM6OAioA3/PRP
f3uukt39uuBf/ARtGyqsuhdVUV2QZqR1AzPV4oPLUErSJpAG59/MbPuuSBBGxusVzLX/GFZqa18l
Ma2lNQmJyWzq9Cd8wwyeoYI+Ca2OtJm2Dl926rZLK0z9ttzCVOUiO4SKlTYyrcPfNwMietNYIGId
ATmccB1Pj6fBASrgOjZhJ0SLLlAKvWTtb+mDzwgpUQR1N19kITSGwZ31me36V69jQEc29pSwYPex
OH5RWl6sqI1SnamT6PVSIf8zvE6pUvOFc1LoftY/Jl6JPnmqh7MIz2k6WuMEK4yKjPuGqLeMDEMl
zRQmxZyL44IwtXmV7EEFE7eKEHaK9wlmJChKugZ5qgI3iHOg2MP4ADzJZq01iMMr/DwS2aPQzU19
8UEaBxrjDyxyuG+NK9C1sPDyC6JkaCxfpE76znj+uRpYlVd7K4TXqrHAX65mq7outMBB5odZL2oZ
TzUqpS1QvxFQReZlHhjM98TBlEUZMV4jVm4aqVtk3teuAUIDqpj9JMfNOYT3obefcvP0N7+fWuKH
bcO7lNa52x93KB1LUpF29sAlYfb4rAZu5MclP6Gk47Vw4+A87/eV9xZdY+fuJtE0rsscVPJ06T3f
vX2OZzt4s9WDST5k1o/SsmlK6O7CpP0OFJNWECm9li4+GQKpEjdYVku/UxK84j1nHes+DJhPh3IA
GWczF5CeWBIbNqHtH+Dsz6DRJMFsADahKF18r1CgystAfHF3MWAVw9VONPZn5lt8cJJOuVeQc2pC
oNQX+Ut+NbKJFD6Dec/1/fnknlrN0OkNn9/TL0uuqAxJLCAEgw3y/9JCM0MNnUwF1vXeHseo9uMt
rI3ietcAtaJG/pdhRGQK9mvjXVrbOHIpsqW5v97hrpKELg3wcjzVdo9t0ptHOcjE9yW3Z1gZwbEU
co8O2AbYRDdqGwNYMQaXcH9p7KwzvIgViPl7fguTi1b5AbB/7AZxPzPlLiM6Pei6IQQB2heKvdu7
DWIg6bIKRJD9MgJhkkST2AjMPj1uC7oU3OdRpxl5XERJaRHDla2x7V7ukjgcuKU41f/tWEM9wNpd
Rl6WkxP6gdimtXmZDD2bTKHvJo5xoEs4SlLD4g70iYf/mkS7r0stFzP0/zsZ9MhiqWDhvb0cVJTL
xD2bmpVZTcnPtUZfSXkD32ZZZdG7W0/8kYDpA4wHEfPd9BNQUakWISh/gaDgvcJzJEDtk8OMzcZE
Z5BHr57P9woD16gV6+BfCo0vMbk4Ex0RH7ZtBg9k5wdy/2q8HQHsXYDrU5fMyeoftRc72OmUoGRv
iAOd6CT+WSFVp144fenAXQbuvColfR4oLdGlcooT6vDKYGpiefvKndlUb2AeW6+BKttXILzBVNJC
mOXMvUAEFcbhFNMLySklYa52zghx2msjqz0NYKPb3h9RCwj2IK4a9tjSy4ar6pMGGCQuFSgePxtY
E9tthH8OIfVIst+oUMMvSA16LwpB0F3z9rzPZ6MK6qS0B4zQUqyrnHDGT3Jhj3i6i8yAteXZZuDX
RpCME+X6Lb7RtCPFmRRDrj5CPfJ7K74GxF9rEGWbv8vdfjz3hNoCDGoM933ShxESdB/MM8mgPJz2
T3eKUPvJvc9WfKHFbSl8inM2CRETkttRE62YP3aDD1/eKQNhBhWKCzgxXBaPq+ya4KcSTiEO60YF
xGDJA6fzlNmih/awKMbtkT3AoiHr4tbJtJiTMsBEaMb1PuZ/joRIZoSIbY9ezaA6muRQlhngkJv1
4H5Tof3biy0WBryZVwc+e2dmNgXPRCgg1n83IGHddAbyRp0yX4JxsG0juXcNY53dGnRmg0DCoXLa
cdunkhvCXjXV8jYuy3BYmx8TIC8BIDJLO023/VTPrYonLbgoJjyOByzqs0suPKt8Hi2R5KFVEkg5
SAD9hs0IKtR/ADZ5vII+OjeCK/sTbUaqDqrhf7nj080C9PrDNDsJea1MNqhH9g653JMUc2tJkdQp
T1xlZPYBleyJK3J7758x/+rOTEKRfSGPMqDyVLDrfXgHn5J0d0hdaaz6BK2JuP+hDrSz2E4MRhYr
aAJiHIk3zkG1KC3USKZvjxJDSHtK/RBrnrdFKEWhmG+M3LGg/LrVoTcq/r+PEAm2bj97iXUZrvk+
EQLF9lbgQ+KFV0EkHyz/d9UyDRgJYW1fg2EuTcIP+XdTEe7WqksMfUm7F9yj7y3Q7SavrFvaeQVw
FohS1JgYhI4Fcv+w4pL46UEPoPbBBBO1E9l5jgVDjWeR6TMt6nZgNTas/mAaq10sA/EBJYxWRn/A
xrZDL6/Lnay/C9fAgE4+YrIzHMe26FDcDKiYONVphdIPMcP2owAPpQGEj9gerfW/7PSLXN58BvM4
Y4ocIjE9CzZZQ8YkCrxcyDF5sAyWCd9gF7LIRZH/UnqmdOCnQR99xooOUulC0kjlWlQQVjUGmuqb
yxzJxNa5GVxhm+LemoAGGS22TAFC8NsqxDh4OnMx2hfk7ugtIJdfC3KR8ydwnujCmZKe7Kodzoec
B0utyO8Xvgm41KghsZlJmlxHReE/Og9A7yeHwG7AD8foOCD2r0Fs+Oj21p66VpBllDcXBA2NqnnG
NWe2I38Rk+oX+dflF4DbgNt2sd9osxaPFSwIU30IdwswwEhKHw8NAvnrj8HBGDtT2Jw5q2cJnbFH
63oKV5g5XxavNYB5u4EswzDY3qGs8F1Fm06zRLXkXB3cQxPPghQMVSwtt1c6J9YHgAVKl2QyQeeJ
EkhvmA08c/gMtx4CmflNw54PrtTWpdP5o8kt/C30eJ7q4gMCsfS9bZEBhiFgWs2drIkZr5xn90wN
BV+pIfrvROnUx88OryC31N/gepPGgyQwrC5ompc3Jf9donTXRob0uh/Qhi1hQaaNriXUAWRBJAD4
PVAORz0WzbndgaQ3mPnvgscffKlb6FiG3DTW0q665RPHcrgKLilURsZx5AulTZ7cG4mMIkXKSe0l
WCUZ1rZiBNyZempN46Siyqj7zA2sVxCeaXWSDdDu1HmlrSYA/KiDviPL4O+z0jzOyJRw9w6qxTP0
GLYk/NDkk1SvAlYcLl1TRPzw11NTh4ODWId5WcQveaxnMzrn1zyDFvp4gkxNTnyqER8MmIOM97IF
6jbdSQvgDu0bH+dYbdhYzqN8GMon/hPrtB/VUhJZTuo/pQGkCAhvt3wISOLT9+PMJGZghIK/vMc7
w3rraxXZb/sX7DchmCOAfj4OAmfXTeM+i8wIevm8wMdN8hzMTQRrfartcGbmXnzevYfdvpdVgL+4
4AN/E4eebMOxGmRL9Xmo8nB713ibVv/mTrScUcVKgNe30cZQ4krir7sZIDy4kWhRpRH/UdO8hYYB
NvMezvyPcXjuFQpiQJO+mkwbGUZR5ejxUa7PA4+COHFROPRX8MF3vryHmSyPPc2k5BF/rJ/TqeEe
NqWewZ2VUhbxHJXNFgzD/NT2GPoJqpMI2P+eKtw8XInqjQOoPui8vCuUONWc8u/RbU1nptTrVXhh
fSAt20f43DL+xhG92h3qqgL92OJkv9w3ILbyg9bixExG1y5kVL3faBEB6dOYb0/LMVG06CK/qTxq
cMJt5+WK6JIaAlunK8rAKLQonHJXssJHV/NuzD42JMiRfYXj9y4aciVL28HXOR27UpzB5haZwiC7
46cLxmoZVCaYGKi2BVQ6kzPX10vJAGhgV8tySM13DVQnGa8EanB8EKXYftRLj+zIV/R4tOMmenKb
GZCHqj5m5k2HVhM+spDxS0tKnssPjzFU+oT7TkXRrCCPyb6subJz6Wks60aRpvaD+PuYuecYBfII
u9B6AHoS4+lGs4cBjoIDCIdV0M+cUn/vHJlUNRbAIzrOlgAj5GtoAdwjWRQoU/nHgMJT+MaIXqU0
GiYoiiAYVyCuU16PR/lC10RC5h4GbFk4wrxYjO7sdc6e1owcJeB253/fsOCHM+pRSDIDJfNS7/XJ
pl8LtFPg3xx5Dc44Wp6UFKy4gqykoo/ywr3I3nLbezFdt2gg3Xv864/t1XFfBpCoZduPrgS/n2k4
BV3vHSo5fhQvO928rHZ8liT6I8KuVpbYUCcylkti46ohV66FANZbhuqswLbrakfFGNxDivU5J6PT
vU/MFDMG3/flvC7JfIz+yErNtFIdRgs4ZMLxIEq1Vyze7cBcoA0olxKtFELSBG15uzhMa+rZFDyT
Ni5ciIBZ6zSTmLIfn3HnotQV9k2a7ErOEvdVV4ILbKtcsSHUIBtYcNLM1QXL0WSsdvGwrVgTddpP
I5tzY4m6S7lAHukBKyFL7eU8v207b3RTCKNkiiDIIa848yqVr0gxcb0+X8opPPY0o2emQWI1RXUE
sOTGlzxaZZgy+4z1MnClqzm1IDcpAA8/mEJiwns8ctuC62zdgMM5P2Fx0gkjhOnNhYKFepfgcR1a
0lhkeNjs8eJYcgliMfRwJcLWNlsTj7JMLNn9uITOV/Ll9xdVlOK1BmEbdrDhOiRkqFLUUE5NIgoe
zK4CeTcUJ8GsFuTy+hJwSn/6bsDK6l48goVRRyt/C7GzwRsOZXUcO4HUOqqpprgj1TTR6S9Blwm3
RFp4jvO3synuXapYkZJANW4alm7yVO7zUiQuInqiB+mFHGZd+p57F9qTWd7Dp8YRPhsam/ubXFGh
biff9xM3isQaSpSxvk1XJo7SRlWrqSuPVxQYTkMt3Fp4EegJzPMKeSd3WoMqlZDyCmzIbDwBpxUz
OZtGaTSMtvcg0sCDxRVAFwQgZ6jlmYoNPhvx9v6A6qYCUGre7kkMtQVzTnB0so6bP8YdpXCv8Rj7
VgwTr+XEq1h886vsjsA+qMIEMZ8t8Eqy4zcB5HhILjx/1/sEn4oeb901t0fhjRmM7ybszyJ4JKVl
u7XlespUtgEGWljx6luKJIluUDvMJqmJYhS3NwYQtKx/n94R76nAfIaW5MeJABVXJZApmKEqU6l1
87Qu2NvyiUQxLZBD0YhB7jDrQ14w5D7i4MZKXW+eGK7/6O9sl4wA05dRP4ugLAmCT0QvoGg+IOya
vrUVwTy/oY39xYkBHJJjdTkx6C052Iwhir77X1BqlAxRBpRzyP9H0nID0AYOD4t+tPhqeJQY5YrL
R9DDP8oNFCq9QbNPAY9e8RMxsgo7GK+eMuTdr00TjNSYuUI3ERDI9n4nUu1s0bftEFIXBWXnJoFo
4lUgGxMJsQpnyNgrnCwzC4578Rv0ZiaEsg7rHPlzlWcWe3ERtVj6MGYk3+vvktpvgdJWUERVYJ1z
sdMiv5gda4tZ1jodJJ+DRY2L0/UMc0LSTSpqF56teyrsiP0ihEgSHWHAJHVtSQ63k5/X2T5aR3gm
huKf9Twux8jpohMG4pwbDoS2WtBtolTH3k82BIE9tARX9s/Xz6CEFmWeE0yek6UNTtdUGnVF3ZOE
0I4xtk0RXRufN621/hD1wcDzFiXjT+yb/dQOkGq7ofykng7UBIjNbkupMUP4RRfi5iDp30VIMHdA
Md1BTlOFUoMOaqe2TnADdJ7Qx8+gXbNpcDunTVA1fkacVmcA+v1tLh00Nd9pfx7eTR1sQYFrJ4Ic
6xXdfAbs+QLW/j5pDcG/nFbD7zpiaU/5+kVtlXIjkDBXzvKWZGx9Tvn6Z81buaE6m44uMv20cwYu
LfPu3vVi90LFe2cUYlRtNY8NZPhcorxyjpha9831Fc7H+bv/knDUxnUYJ0SVXxlITlKBGjxdZ5ZT
/Ak4joliPpikrlpbqEYa0Mgbm4Z/ickbEKvmCL4tTuVx6DCFyGDisQn5djK5UCHb6NhRM1zSbvni
HhTy3aCOoyQsL2dGuSRYZb48Dl6Yk4N/mOX82P/rABIe9omIXuU9A/Zs9n/4ZhrMi/Cfhf+fD+iS
mZY/7DIG4zbBzoAUoY5UMDNCg1iw+gjxp3jE+RumHqbNL3AbtIQ/uzOFguPmbrXrHYZUwqVtgRfz
ZHM568mZZ9At7hatYsgwRsUBszRab/ocg0HA9JNmJzOGsrb3YtVVy27YXXfWj74N4q4Dgs5j7FAr
rdg/dM1aboWrs+R7gNs4Lm0yHk/VtNFrf/ddreqFhbjIwj4JampjtADh781wbOXQ//qCiKVcVFsc
XsAA7ZPqv42KK2sLEgmxD7O/H2XZivCCVgpdB9AvKJsu8NfJIc3GX2aj6XyevDDC8nzOZpkx032N
50YWbWymx40t7eWyPINha94T48B3OBOkqLgImRTVzSJPBmiqgTkWCnnxfb3FcdUEPh+fUlr15J9W
wrhNrrZp/JDX37VODZUGHBj2oYmfLCq6yy5DJtUX4tTj5TldrB2HsgDQVFnq/hhgjXeeJpkk2uqG
f4hmEJZq6wjSt2DdGH+anVUEjL2oxmtDfyKkaq2eYzla2mqt/7OPs9x4z06DCpLM7lN9oGUoVpP/
9WhkFevH5BKnumLxC9PLqmQi4rHZ7T4Wr059Qw5GQGnxK3IZBnbo0oXM7ZzkFCb4pwOMm/rKQL0e
PoQOJtCV7wdS1b5/nGUi1hLWZ/HrfdF6KnWasDX2vA+KObpou6g8YlTVqkItmg/j8nCAIweUV57A
7/U2h1VFZ9dBdjBb99pJpWulfQCai/94O3apt3f/MJMEXm3AAaNgH/ksrwXDQQqkcV2Ry18dazDB
d7NbqR3Qf4jiPLT5OmFLTEZOND93bqp/zcxYN46wVqktlpkkLxFeGPoW5GNniMLQiG4c1m2h2pxu
k27q4l9fIQy8yoadTKEQtS+DS3VzdpBBMD8SgYcFPv+14Gt4eQrZaubcoRMc74rBAI43LrBbtWTX
ql2174Fr8g86Ybl+mWiumZErwGJS05Zwt60atxDKOamXS+YDrdCulYA8eoPjmlPO+2c+vLCBf+IS
yuNOYspBo+ogQ9MMKYVGY29RewPFsN5tw6fsQqBqdUSjvCm6yDKCl85WI8bie6ZMcH3zPyUjHG3T
EAixxeU7sqrd1hsGgIs6C98KjYnKMANbNrQvgW2Q5bu3rZeYfbe7cwZ6p2vnCTNgDAo5ON3t6aEL
Qv26vXhKhGdH6CSPvubCA90lWxlANvTnprP70gSnl3gGjdBA6LJYunGXzJMCKtwjMMvqqI7En9nW
dd4z0A7g56PJT4dt4cdT2eEscuMDZsKWtmykwnuJLW0Q8+rHjxok8N6TGZpeAqVx9NlUFg8Cte4Q
rJDhSTtUmf8H0XgviiplcyVJt3lbnFe4yRggeFT3SkR98l+XOhz8yFVptKtriLv8tz3ojd1MlxA0
pPSBahQCF3EyngiK6VIg75Deyj0cobHC7GR2MOQ3b0wrBn6HqTJiqR85jVtpilp/mCzw1E6ThMXQ
rbSZtYWMU6P3XzxekeNR0hLUV401foalSN0HKbm5vixnHto/rDmiiYl63msNvPT9QO3rCp/FkkA1
weg64r6VAFPoqD4H7oQaflxhbUCCmXFY0cozRtS60i4G871Rx3lF3pdXgbyxv/sbGFTA/SaJrVvA
3XZVBso7+suMJFGszKzMeh2gdwyA5wscJbjtkdnq1E3UruOj7eBcKLdnMiqzPf5DWcqT8F0oY1nr
ThMifbhyzoCiKNA1eqaPy0JVce9eV5vBwRfxrVKla0JYoXMlja8QUyGaxWV7Fl7h88r0VMjGq2sp
M17We3OWBuvT/Vsx/wGZ5mEBq52Yg7qraGVL76kl6Exgt0gnU1Pqhxd9W2+XOJupvbc3BgcqojIe
Dr36UqOpm0imIaWVWyDzTkviNvWO6EY+Hf70c2yKBd3GFs7do8HMbAMTdJpkVex9AqKB98MrXvdD
MQ4oiog9n4GTkPUimsBxATfLxo1HdfEfSvpOCqxL2everkgaAgn5SfAh9ItcyMqKjrFizWHmE7qf
OYOyYGBLYRSY8F2wsU19c6GxZOsbML87d9nzW0efJbUDFWrcWRfpiflJx3f3y9+ONeGtnTuqeF27
6fKnM6hB2BwNy4PlZE0ZkqVlJ9SSfqGpM6raefjscJRs58sp1CD56EGZ1xCdX5KFAaE/N3Jmfupo
eYR5nxGJol92ZiskavPH9wiTmPzKGKqulQQoZtXDIOWX+lF/DHMxqzq5QirDfarlWSJCShlaykQY
e7lyMpMLfNDQXOW7jk1mI0uWUNtdiChw9gEGL1RfIJ/TANb0PeoH6UzCV38cSE7S/B0q+r8i30aG
yS+6pa769AhP4w3z2PA8p1j8fUiaqohnemRA84qJSGE/Fcu9l97Vhs92l7JP6H2Qz3MrpteHrQ2s
ueBwIit9C04P5ZZ6NkA1JjwdDFMwtZI4Txe/hplIXYg8Zme9EFu665AZvwnzz2A3Q21UbgKJnR2U
xadMSjQuaoOYtW2eMod4j3iElhd4jwH5tTD42Jcvpw76i4/elnAVLoB9J5Arf65p0pl6oaNOwEHb
2MaIEO8pAnhKHgKYsSWtwIvfhWQi3dOJVF7vr2mEwNxwOWoZByYOjnq8fQoi8kyOEclV+BskX9Hr
r/c/2GLRFtx2NwXuadMwnAAm96Yqi4LPu9HIOY3r6K8GYBHOvkkeMERb27W43cGEZU3kOOC1ya5V
12XHZnUkZiTABSzdU+JcNzPUn2Mqzkt7Aj92sHBfhmDZuQZh67AdC4/erRa/eHF4XTwzPTQgeSYX
AF/EcCWD6TbkWxYE9EZYL2zQtsRWxJVQ1kfgs9DL4tMGSYM7jk1n57Z9uNQNRKMXjrGtozd51ST9
w+AZQwNFKPLYomM01LRFNT3HpfDm9rkqxeNm7sLiZocgkSYupJe95MdnoOLPc7C4nfJM6IaIa8mr
+2f36NiIQ9xp1VgsggO7xhrq8w/2tyA3q8o/7MiaCx6mj8LIPKHvMKIE9MwghyMIsz2iieSd44rJ
vsJ1VcN79We+2KvCPvJV0NRxtn9NT09FKAwBDomQOQre2kaZwC7V9yeBLkifP6GO0mcjlr+hwkkc
PgWSao0BhqBbfURrLBXdC7fWFMT/JrinM9WXoUnPS1gyAVaUPB+QpqQlPiJIABekZpsqZqQes1Bb
1u8+YaK407/dqM8/ZZiB1q3m72PiZCigmx7f5N3bXTrxFb+ELDNbCBDsNVCW9kmmSS5X6yV8VqM2
yz2JS3rrozGuSaFzCYsPHkSO6K5HRWQzKZ0GEddLPP5+JDhhxUGBJenOdv8Bxb5kUI8eihLi2VxT
eGvqcuH+zqk0dLOjFIyRTye36T74xFP/s4vufG8I5KvaUpMXcSwU/QDRxtBuC8xqC5I1Ihw9Xv0K
h6TbpNVQKjM/jOVYgyLItQIAiRPORbJixJraoo2bKMvaoTH0mdBO5HMI7+1cFlU2aDylbzOVQ9dR
2nUA8ydU+VHDFZbFBFbMOnrnJd83QS/AxtniuWyK3jnOqWINtUzru+sQ16RG4Kez+OMGEpfG77Oy
utgTsSunKEhFgnwXoXF7qodolMR2IkfZMxp5HKDEXe62SBjXsDhBFAGSJ2cI3rhbNj35zZE0qSNn
GvyZG0Ui0GsUmb1qutQPQ3p7rpxT9luOX4u9jl+yTqzZsdsZJ0iXlisbFSihu4rEI5bkHfvZHwBm
GmEGZlMXr7RuXbsprPn1z1qqk4b+HXucmLgGjyHC6KBVxSxZJon8DmFYKpCP1By8CxoNZkCgkX3G
8MuDIQyn+SJis+F4ohQce8WWHK7BzASrVWjYwzDMb5MD9aEdbKRUtTB7YNT/blk78yVYLGJft86/
SBdlVqM1cIklg6d1QaVoBBYp3ZcL+Ky2ixSqBTe3i+OWrFYO8Nd0bRmbZgZlFjkh9jLj3RJFbTLk
PmvYYvbKITVpJYNq2/yLis3ZUM2351cUNOuRYHoe0uqXTvBSnHy/IATl6r8mKNOwApNvM3a2imIu
7XIfeBgvF6wk/3XpyG1oriz6FskRlAZ/k/l20c/C+Q5RkVoF6r13jXkgVEw3V6gGWirosu27amN1
hW8gu5HKhD6kw6bMAx7r76v4/JAXWUjZJaH8vJLsuTSm/J9NCocZs/UtzWf6fT9l9pz56LV/NE/2
hdI2kRctQWGLbIV/0v9o2q1rIG/z8DOkI79SHgAV7pWAXuV69iFqM8AtvjnyeHYnl5jVCSfwd+gU
tyNIw204yNduUSx9TqbAH8FaYOJOzyLsOt2w6xFaZABh0diRbFe8Ta2M2yHH80aFZwojDKjRwMsu
ydRhM+zFKVZ/51ckjoq9/YSN0Li0Ao7yjhYQe6MwSmHo3bMRuAmMCraOs6V4NOzwBXTPYKOocW9b
dCCb3Olz/ov4tQovJZMdW9/N3AyofhoiIgq7V2WUMltVUYiv5bqZilCxuOSDNqxKyaRIkEI2Qntx
E1Kk2WungwpDdzGNcefUflnbmwUW/OYh6Wiik+yy6zJPACwyNHh0yd61Wvk52QXT1ZMczltKZ4I9
Hjl5avjnBbw7y19R7k/XnsfptHlZhhJZHTM5cj6nYN924b8lCWi/iYVRBMdCzuB4Tci8Hsgho2Aq
3pD8L/VIqG8PsecGzGADF7YuB8OU2B3W7b+WsQcub5zaaQ2bkSfl9fXtQpnmzLsvYSvbnIAufEfH
GJnRGDaCy3fHwOdFLgBK5A2iSKqoxiHOxVYnZkJ3nXmQhVgrbWZa1Ygv6W1Fi3Bh8+5/HXADhUVE
sB/ef3uQM6glA7jgjmKY1mz0KINQZF5SSbaMoBuBddEpO61JL8ndULJSBIKeTsBhw/gLq8Y08cV1
WjgftSLrLugvXqkJvfndu1m+PrhutXBnLSCYXihHX6oS6lyRu4oiWCp/WybP/Nr5Lfoau+CqW5zV
kXRo3aSM/l1G0I2V3zoUF9KVv7OSMBvdHFwmuXr58/p1WlleOWzxRrAjmsB+bBQBfPdT/aJdQTdT
Hcu7cSGbpuniDZ9Kq3LshSjHl6RKX5rt9fK/IL/JxGsXu09g4p1bpEPvj4oM9IrhQ9tllFVrm83h
NpyqYea4Ylzj68bJYwXFK9a6h8g7MC492a+YOki4wtQVG+dYjsyqKLUOxPCRu4ad+Ymg0rOCFQ4o
PqYjqlF/V1A1pY1s4Q5nzb3jg2M13wtduL5pN1rxweV+Uht4747tJ7NsVhI2KK0QqyqIjN2xQrxk
XP6L+0dGPqtjeVhr6Q5+Io6yWhxsUey5YFQeU8pYfypIdrYhBtyGw4l3LCttbxW2/544gHgZS277
Z8mylTeTgAblKnQVPftL4i0r3SRzHfueIgd0kmn7vfxtx6COLKGEMum24s6CuAfQpl+j38K/Bqh/
DE1SJ5uTxbY4VxXlVqm7wjwL3eHoABsZLJWASlBD+CAcRMTpCKsTcJct67EhDojBgeEyoX4/GIOq
mkgrTptOd9VCxOiWXxHCyi+wGyl16fcdPLRvp9Ewz/3ua+nLvn72MjA8JBiar7DONAQG/QZGZdxN
NnA3rsMYhd8unR0GcEfcWKAETLwGdF29NaBLFwxYLouDmZAb/Un3rKf2xKpOmu7pgjalehDcnvuV
2pWe11YVB32TDcHmxJIF5Jd7Xv4csm2QF6j9XKZn9WsCP3eRbl1CJxP9paR3/FblVh2Pud4uPI54
WbvxYJQnYhgQCRq0CnoO1sz3bPzJxwxoTgK7DLn45l5ojXn349qqXRRv65cDFPCsK03sjEU9L/5K
1/eZF5ccv3MLTHUC5oZdRDj1iTH7PrSBvgcueYebmsE4/8EdkgZOuJD07xIRXITVMQ6dKlAoJeEK
pd359vm+8VorH44HLoq8Hz7pogfAH7t1o6yo7Rr96VNOejddULrLfazzNeJaseRQ7S1gPUnWWilG
8G05miJaP1oX0kL160/rGXNDkYxODKCpG/wV4Bkh0/4OotseR8SAB2rq28aMM3iWKFv1ELioI1bw
waMdKJcpbcld807YlCAiQSEad/h6DtjkuPk+CfRBc3qz887tBhytN0tah9fktjdnqz1XYGZ7Tjy7
gAHXgWV2njMO1MDf9WOGnT1gSemaGEg2P1kJ8mMAN/njDgGpJvIKaiyjaDrLpxDkKNR80IsaY+6n
brFHacRCqhQrOgpRqEMSFQEFbdWZXvGOggmDJqa/pu3ZzctLSMdJGrU4IJv8jhmV2zYRkAC843J5
nwKOVkLk3zZfq1m/5tfbrcCZTMtDSrmT/gCF+SG0hGxbX6je+zdT1hKlFeqocdJwlP7P18EgdE1N
fU7kep2OoXTweKx5ZLY3srrKvNpHDTPje0i44K6M6lXjw5J9eR/cWncM9RPwMrgf7l2CyJE/k9mG
9cMkUo+Cpg2pl+mVc5dDG26pWZpD9l1y440SG9jpLYVez6HzDLWG7BpTsiTVVzoA+WhojdrXrh28
VCLGAVBlOr1kezXKTwS0FIjARB5shNCWXtsn5Q/mFeLR1YhSgK8JMPzfy+O0+xa5Z9D5v1j29eli
bVmIWjeQGg0ShB78ia4SaO5yUh+WmK8N9gaEd7Bwwz+iUOn+byMp8waEcvpkT+W0TJb+n5Fjd1LZ
pCau8QQA1pcdFDDnReGp+KYTntovSCD488egu7OAZXtWCWXROdn5ZE0bPpv3k3Yn0TFdv3Bj5bXq
9AZ5gyDanOEMPr8iOmS8YVWkUE596/ccV9oKrY4MVE+mw0OP2VB6F7kLwBdu5wa3xf3zv1xmrOKl
GZcsMj/IBncwO0JAKahdp6DsQeIP/HBwUQWejnS2Rmx2IywFWYKM94ok6roAY/wK8fqO11jL9onz
5Yk2B9hb3j5pbkoMmBaU/q/Ll3+F5CHi6UygVxk5w1Ivr8hYOTpKfTkhGSS/s3qku9nLBxvbRkYQ
qvO6BAnTRa7/dR3AtsvE6W5xtuuI+tN6R2Txkwa5mTFOrqCQPhO1YyHg9B1lski+uUeGUZL1G6rC
K2xf9swS3lYwkjfIf3OI0k4L1Fl+e7LMdvtuPUxjK34OWLKHaJ3Q6ILJQPRWfi4g4/YVMgG4Y2v8
LVjXumJGBQwLoZsw15qunzHh7kRuS/SobrzZDH/2YzUMCqHfi+4MTUukVJDkCGEK/yAuXbucChMG
TJE5bj0v+aBkGkxJhtJ6i3+q649yNAXdOlhHvsvJT7nF2pnWNIDS6AdbjTzysmfaJReP7+4X7hBN
Wu0IEPKykBUixm1d0O8cD5gvjPeWslNoIm6YHq4sXU9wGpp/8ie8JxV9McMrknqtc77qO3gadztH
VwT5cuFviwu0i8J0Z6Ra/L2u1wI2HiQukXz4+1lFox8LPy4kE5B/59OV380OXs9uxdc+HCMqOYCi
Z37O/G8HtdHyeMazggG5XnrDApqGvhk1hA6XTRYlhAifOoPIDdpEPFY2y+754CMozpEFrA2GNtod
Lbwv4yQg+JLBEISLturWFYt8zqLvTdTnnNijd16eks9dtOR52HFNYaTrbNOgXQWm/qxv5YsavQwc
H93R2fP9M3DaAE+cre95DZ5LZsw/1ur0rBPGm4dmJq7JR33WsHQuK9Hb4/1Kv3ArimstZ9Nr2q0R
O+TNFT7EV213nn8myZiLyMhKrROx41RMRAtLeKuYQS0KIzVgmhQpRICpcMOKAKFvktDT1GTN0ecS
iTmaL1eOZvwKiX6PfrATg9KowVOTLi3pch70WAJ8IqUOZvARc9r4+BLbcD6kvoFTcAlQWZDw/uYY
j1Wm6GqlWLeZ3prALIf7KCfF5ICZ2Br+b83eouYdnUcRG8bNJ2KmfN8muP7Zv42B+PvjZQ4z4hPl
kRaDobrRIGqtHT+ovq30CS3dybF/qfBYs7UdRaaBvYUk63YNQQmGm/aefGdsbGUh3SUFCjqM4ggK
z9JguW+B6O2pop6mffpjisVjpuwhfwLdPRhNjsMc4YwHbex0h9bZs8N8ZlntjKiBNMweCSUMnTLn
JwezoUdSjwpK3T7D4tmYB/o/kiGt4JnD2DWe5y0vPZyqAWv4xBefObg8mBNSATsZRa9sKizqVbWB
Dmi5lKStPmbD8PWjX+2PAz44mfo/F4CXyCdpGMYVaXrSHB4fDlKuwc08WJXIBsX3Xk8Dn7aoNUF8
II+ZSvLHhihm/ouzt15vOfGgPJeQIFR3SvU8xorhZxNDQG+aAvwM9HQpUsHLIW+fySFvEf/RLJKn
ohNIEO+h8/+O1lXhuCCGmSSpiwRNxiZdnMh5LZB5Jpm0VVCz2bOYOTt8fwjukxpBBqBrTfBzft8J
lZLB3oQ3FllzQXlusEejjdgJ6zjVw2T+GQTDoT8ICdWkBRoCRYGU+RKh3TbSrXp0pemmQ3OVXVk/
ZN/mzSW39F+HxJwgwlcREVAdonPNBuKKtRcJQ4xf+9Svf0J7mNn5JGoj6TM+1XhEMzFTIkIT3Jas
jhGEgTcfVzxv23yh5X41195+MzUJ5GtAsbqxR9m+r/UKoiZJ3mDWqzXTffXaCrzBDfTgDugNkuXf
0CQWybiCGM8hici+aDzbnVdg0fOVdKC8ZqmAbpvzY9pVxQc3myH9Li/lK4MWHbVdJnnshOqivHgK
y2GCG20zsJ6UmfCOe0sE9ADfQFXqMUrIDeZmi311AdAF0ZV2k4c4TwVetqv5h9/FC/5SZW27cefP
/ZurGGbkOjip7x2eLv/L/sQGiwlb00ONYpFm0/UKhGykr0umzxeBFvt8M0twHj9y3kV0CDvvCOQk
oOllm8f1jS9PWlg5mbunNYl1/BzhyA3naBpfi1fUaGvhgFgSV+o8NwDTD2Y9c+EDU9UFW6BBCzBs
E48yfx0it6+1KF6Bz+jW7JxU1X9LJpAWIAbA6qsM4klS9zJPdqn7T+9ld6INzKuWR753bPeRlFtZ
DhfSDbXotaEs7L7wlxk2xGe6Qzg2oBeHtsQgCNgXhpfJG3Ovp2h4EpULs5RJvXnEjZD7wDD/mYcD
jsb36LWKKXzSAd5/YmIEeKr55kJfBKENEEiW6AoLgA/LC7AbkplkECw7bHclsKGGPdOo4YalkgZo
qfB7msr1N9o2NXQdw0g0mTYYgM5Aa1OmZgJJ3/ssXKnuUPUSTow/rpjv8Q/LE0l4xqBo0gJd4xlX
OIFcttL6/4cw/pVyt1VcmxySwzQY8i4Q21plHeSpEKfgObNvdTpC67IQaAJ4Tw6oLE3JB8WLQ433
EThh4KCxXREOxMoDxgKQlJLgci8Y3h0W2eruqFfvUiKwxnuLD5p6+25YLa8YnpP+ZhYcQmJeXUIa
5RWhM5MOauzMLRj/mVdUGiKPEmqyAvxHXXZVfHENSASbsPJKA0kA2zNgZXpb1Yj7p9Yo8VvpwTQ8
m3BKmWVeVhbYTW8n1Du4wBnZ0tbjyl8fIe6xDyTsE0ARD6nhMTLykLnzb/bt2r0ODVLJS1biQCWb
ObFJMz0hAE6JP2W/L/hGju6EFd6RSIbmJ+6jhpUC0ZszhFy1/hco7rzNxAX1p/7wmE42qriZQlIY
qdXTBGhkLwthd0o1nehibvhNBWoBeLDazWPNxhGOQTV/WJ80Zt9warRrZ+iha9RE0QhyYltG+Bu+
BIW+PJMbDn8pL4fZqDycqEjfqr9DX1+X+aTWIuKgvD9MM5B5XKvoP7MhrnoVsIAB3xT8CrN/9IQ+
eaj/KX5wAZXcSRpJrSe/8oqbzK7Mx1ZUXpvqHpVlKPLVpkpYUQVL32a2bnwDb/2KFg7p2zDpPdgn
zCEHvrlXeWBackTTnoktEzc/rtvw5Vqw/00s/8GuPxsE7XSVjuQAzkjdoARivuBZjPVE1EDIZkiF
f5nigFyVWyxnUF+oKh0mubKjgsTf4iXhKlZS8Io2wqGrHnp/23b2aNjwDYNaij3mgdl8GmK1dndE
odZVEVPDnapQ5pwOYrNkcnUd12yFUPUIpnTo70O/4K0yZfnv01Z2HOG95Ps7QimuXFKvVhmk+XEP
ILmP1k95y8QAwyl9U3R78KGIQPVKAIIrJW+bZOWVKjCEGptV2Xm0qUxacB3Xz/YATcd/rse5UeLK
bUxeVu7mNRh2GkY2FP/bx/QgAGahbdrwwfgAu7GJQ9WIfQJUEjX/42zmszU7ob+e5FuxUipIEWBB
A6exTAn2lqAVxlRUziefMOwXUc8Im3PbznrL0lKt3u8b6NwgOL69R8HPPhWhrVolyXw03LLtEAfY
KX+dTa6f5J8GNhZEt1AE+5jLVS2cWI8tcUfFeTuXE2kAjlqo5Wiz4gCDNrAN3BNA3LoiexAKHt3p
YsxeQHAya+/4Sp+W5RPUu3MCu8fCBwRDd1wzVF5zY2KSp5UpsnQNw0weC1YAo7qFEucXUBz5GMrk
pMPPzygJ25M6YFskuDLEqyi0Vnby0iHONBBbnJ/0735pOvZsKnpInLUaXK/I37WCPg+C53kRnH5C
1Txm9UHOnQmiOR1kmq2cEZz7K+pbWTF1rUQ3fmHrs0KKRs1VWpVVM7Vow3puBeYGIWN9WvOExXuP
9b+sQj8ynu7SnWu6Y++xQWEWubzIHCn7GXampHfZwPRSwZKZlZeYmabI1Hc5TbMxHbxDzioPYHdt
nU86c9cqYQVoDJHZw46DInfz07WDKbqPLf11/K3WcyvcSfrnEFzH2sgDIy9vvWQyjFKo0VThTIVX
R5dhJBZGnbd97luX7VxdyUF7xi6IVsuspLTp5lb9UKNLxTyrKvKKayNALdPPKOT9bHBCmn4HgCgx
0GSJoAstYpkewgXr8fZNLr88MV3OVyCO/TqoZfongGa+To7/IqcJvD4lqh1uJst5QrghZzoAUIHo
8H44yWzc2MVpz+0FaoM3rCeUjR5hfA/wruIU2esjwzu4fu/jM5ir01yHd36dUUARbMFsMOO4vz1o
l9zwRnUjF+pcscV5swvyjDlfmIDClQdYOrDR5fBtvnbYkJnwuoVHxjdfXgexGbC/GQcOdr6gS4ob
M1ak5QYku0UOnL0mE/6EVA4weSDFgCWyCHw5evkoeaut80kvXjQslEsxNeUH3ZN5J6FXUpNpmTGK
TBnGaCf48vpZJ+H/ck4fyVbQfhFB14o4es+0paYDE7af4wyor17UwE4q016xfHVXBkLpoOKoG22y
TE1ImJbXph/DkZZ6o67Qp1O8jQ1v6uQT5WscWcfH8Vmj+nrALweeuji2GPB0x7NEeRMc15epxiOk
9kHWsKf2ZCqlsecq2K7e1grIwBVxBlAyVbqravEcpeYTMns1TKKrgA09ke08kn9eONGHyHOh8pAq
MW8NN8mmvcgmYYfbH9xQS6ua6ABFrscyewCy2YGwm6tpIv9peiPQoDu7M5ZjJ+NhePn7fEMqdvF5
6Gtyw2CCiZXpOfhE1OgPjQTf9neuYdFZ/7FhAnrEP5Atsi9B+4mnUGW1hPSVSLTVISjE5amifh/k
mDnk4+9qsFXl7mFx0djsWeE8cbOwyis2FXRbPtt8ZuXJlLbeJc/AoZwqPv3QcW3Bl/FO1q1NFg6e
lCI7fzta1AwyCzU4yt4BqvSAIz46dUNSL2I6/LPGKDbG969bxd+Hv6i+e6V/ZygoLyiCra3JvnfB
aDTHgRs4x06m4F0rtUNN/u9Gd5Cux3EIY8NPvFmo6ZFqZdv8l4n7d2fBo+uGsabPq+dSP05aa4D9
gP8bAyz4URwLwjLPtoCPcpLZiPmH1BOOyo2enSGTJLus8GMf9HZSVKq/RNB9HGPa9lXoDLwX87Pt
X0FnXE1L57r7o/31soumY/BGJ2e3nFXBpy5z0H/hCoQZuUCTNPcR3hVLNZ8XwZqzKr5j51d1FNW8
6ZlQPWC2HkKV9V+XM2EloQh2xo0UEhvlysDAT2P+SFdJzmlkc8KJGBUAxyH/C4M0O4AszrUWstmz
Gn4UeoCBuMTmxu5JY1jA6p9jhLAuNh/rRHUDCpapMSYXYWzHOJCUjoTmp4AMViFOAFNjRlmtqCUr
OyCBA+Q4kxwnKxaA0mbDbs2ejieRmtDJqegvRpRHAaWnvDMrZUikFSyt2mQwq3lOJqo+Oa0p1fVT
Vti5QNieF/HOwnnw2YGcc0IrHOTQ0+pPRZ0o/kCl0QwPUcSq3ix8xk2lJMYpFBqaGMkx/WKh2uOE
PbByyGxuQzkomx1CI6uJ0UgqptmOiHoWlL6kM85zkoU13yduIwcGuR8Be/Qc9iUzuGV29XK1tU/5
YzTr2sRgBe/Ur9MnlJpU3Dt4cLdZL4z65x6ZVid8lL3cRrulIMsc/+ZpNFkSc6Wj8LWUag/GwKBD
N3s+nDRdRlzZI6kNLUxJekrgmcKs5PGuNxdrU93uKkWhF4K/rRJfpWQcY0ksCSQHdRr/TMVXkhuA
1ywTNeqDypgGXh/9SMJFbPeiCmIoiiCFgbXamYxtNwMDLNzSLzNzxs2mJaVCcUsPW+eT4lP+D9DB
On+FpHSDQDaV9Nsu5CW3KkbCo2wntsApkOy+3AFRaXmiEajSwQb2WNX3NSfKRRTBUTisvBbHq9J9
08hoyIcGs2U6j6hbcNonaly7TDWmbQYa6y0IuJC/6VEsTXaT5FYB63pnsawgQqQoBN42VXVuSzoS
ayIRjM8sVvQNhEFoZX/JR/R47eXCI110fxLmeFXQJR6tnIEy5yG71BGCVigCa/d0lJoTaYZ8Mf0v
GqSwgwzRde20q0GPvOF+RhNGfDi3QJgNIXvxNesgQCzdhJu6r7cf0pvjvyWVTw4ZEHVHUOOFrf5/
Sk0Hz0DBzCN+TiPMh0g2AROecCfg1kdDNyMm7TU5i8+JJZK5K6bCX17ZeMTMqXDmpzlWpCNv5LSL
y1FBwPH51A0RwLfWa8XSm/WCwQ2meNW5pE6GolC9Ao4dgd9mKML4c1l4MeGXt3Z+l5gcq/yCmiJt
oI06Vna8QFsWRBqkRclEYc8AUWX0xl9SSDFc4UXL/4GNyotVE9CvsoC0ywt97GmqGyxx04XaZAFY
MXsK6WiGuhQ7UNfVoFlj8eUG7vhIyOm7qmLHPDyz+iZ36Jt3BKGkzoiMfpdFGSPCtSv//Hue4+zo
P7zS+d128vcsndNoOP/8TxCCplx42Xt1BBof8B0B9aKdJQb2r5imw6h4HMsPTQmbWjBrlqB6Ovcx
r5aXwZRyX8TW0PI6S8Wx7buc3tsoC3fQzEhPjJhGaySCfQmxn3IegouwbJ98qsn2U/KezVyp1AxT
EJuCdagEneHusoz3rDHt0dy7F8rGkugHAbGZEpxm4C2/D4z9c+P0ec1nxgu061YfIDwJnJcpDVsp
3ZHT+wnCs9LLK2bKouPl717w38jaXGyw8AzSdMy/kqZWdxe7W9UnmtCjHZVnO2a4VKMqhx+kICc0
rTkfCkvZTdEKuJ43CJWfh3iS5uhnkW+iEZil0cje4xw60zF/fnFMiOU6aWfcEFJdGxopopNmHP1g
OQBwjRodGCfbJx2CkqnVsYF18c5VMDyEC5QTthLOQBg5mv3YmU9yiM0FT0l4X31iki5gdleVCXvP
+oqgLpb46XbIqs4+L/kN2WavPxYZaACTreSPlzrdfMuylosk46WfMzMS65bTdMj/b/dB5TI7yEc/
aehhQDeAeuResKIJ5LRzZ5UPTznUjjrCagScHsi3ltrwGE2T43y4bqSHA7/2tM+XspD0OfWcs9LV
ADK/9S4YBnptF3uBL1TqsOdccQF58mo4mivqD0KK/SL5kp+JquwdTgh7qYLB0SArJSBbkpfCgc1l
VHNcL6uuLZn8xellmn+DnugzSJ/0R8dHt4ZusWnGqhurCV/BYNbvdFDjDJD/PWZjRgXB+SasiyH2
91phPTO6SNptgXCIn8q+Qm+1NhYQqzXnJwUDmgTbRjnNWEbio9+i6bgJVB6Ukp869ZrOHIVYubqj
q/Cs5M51ydhc8KuK6CMemIbJQ0sxTTNr5bdssKj9h40EyaDSSOQxGVxF4cAVjv4r3t540P804DcO
MBgyZb3p4LoMJLZPT0Bk0L8NzfQrdjaatuoBHBjQU+PJzm5DuF+eG/b/7qtLD/2va1ES782+jXin
Uv+KbmiUcG22/PTRf4GT/sUG/CiZybSBpnSPhAADk4f6QtvoIn92UPTnIeuUAlpj40rp2QzkVpM+
DJvfL84abLAoGNXpw885+7NPg0OpsNANYEQCPMRVDdm4PIEaGsmkMnbTU+wNqawAs6FA1AjX3D/A
mlwfjnS1gOVc4mWJt7F/OjLVrGIA+ERfrxCiggf6aGCM097VR+1B22qZy+e1MJQIB0AVFwU2LNBP
jSl2x/Z59Gv1/qRLxLjgLCt4gXEFOMih70z0jhbNeC6XgcYkESsfDJeuG9VgcsP6KfEtkxippEMc
NK3aGeA/p1THaGOOOj37C8XDAzXAuS5/9AnSfB5IndLj8oTe352wDSs1uf7iXczb9/sqKPyIDQ0o
7hwHodR7lyXvv1tlAEB/p+kzkPqhU/RrXKT45J5ubstjo5yJYNeypyG6AjNPsm6hZDzdSg2feAXT
NsLlB31xsptz+qb6p9jBqSVAfNLPYZ37Bp3ZPTnjhpv4qmqBkQi2m4FFpfbwcpbGlFltZSD3CXZn
MoEsyapesW9mQj3av205OE6exg22oF4Lax38tcrL6y9mK0mCHGl9YP+RMTe8mfdbFd/ty+19Sgwc
BPenxoz3O+w+Smr1UXPpKaVaoIyJ/r7MfFqG1Zmj9MvvUsk9fqVbYnl088gZwqcAsQs5AvZIChsT
An1hxru3IfLEBocTjOBXupf1H0Qv+Uj6yWlUonx6gB08cfXFspUgxbbZ9twqVdUgBXhFqlSvawlA
1WkXDH8ThJlhOfUnl7hz7ySsTjMqira94HFP2oxeV6ZVO8iE3uIZx6MnR3++hy7XqANB2ekrLidM
wuUZuJ0s4ge7lTB+GSnkYtsnjX5KW0tHXTPy0s7i6kPzTYkAUeX//z30J6x+TgA/XkdawSs8HiXo
0WXAY4gwdXyHnJR+D067B9XFxf9xRZAr6F5OLkpqcqnqbactALkAvmDlxIU6AXHpVt3slXphQ4MG
4+CO19KBNLWIA8kG9zv3Mslu1tij6W4A3PGgXmAo9jD0vfQkNyTSV8O8k1PXeoxXIYohpfMLHpIm
YmA3hn561L0iaupiNMkrvfkaLbf6uI+m2qJYRR0kwUNv37WNMfhsIeAgCbFH8W+W/viBLeJdmwD5
BmDoAqJy4379SHlME3TJFfN7r8W5i7Ibuk7KkykitduV0vqcbJAuWiR13lVV9GIqJeoriDm5UW4z
PF5GSCENFd9BYVBiWzDcwQiSzI9HgGOk9J0ZlmX1GZ1n9bRNZtfUbNCOQLQ4WDCHjAIvx+IXhWiB
ZQxi6aepA6NMTjpBiPjXQqhrmUGfqmvmeTaKGslUAD5Rg9IaUQcwDCAlxSojGAI3PMLuf0pknbjZ
JaXLBuXyxicEs9yEibVY++fbXv5TVtMgrhnhEmhjl9aBMzK++P+6/oFJdMWM24yfVrCegTka/Nag
LSx1oKYmc+hfutyXQUxUVRwEF0TuO0WqDwpewlXzwfJRw8J7sBmYLlwbmqK4QxvvYEtM5eIOI88C
o4qmaK0jY/bBk9NPeee60fKyGlc+yHCk14r/SWhItBptSa4MNdLEuZzm+Qm1v+5plHaR3arISVNw
helCFeQVUO258s3fo0YU8n1zsksXP8icKc9fspJUCcTEPpSszSjNchXCyCdsjGeD63KNBI8xCY+C
+rO67HRLlrHJmlgBi1LSOoHbQy6rHeKULUZyaIeP0epVKUF+5NrHjID5LtMtvT0c68EBwh42TgIu
9xxE84AE9EojSJDmdA2wrtQzvYQleMh1T8zRfv8D5ggqKN5z2g/U6/3fo+s4HIQ3WEuRhUePM2Tj
8VtXms7tiCaJQr1eytekNfSS/rBYpYgNOraHcwqpwDEs8KG7FsliuHfTys0t6SIBqGm5d1BivNCR
mbABj9v4jn9EDzROlegC3LF30++UCvrGYbxOvMOU1bovL1hAM9boIE63CCZmIo4rxLAtAH3p/azE
fjSsAxGccWJ5hd0+LEn3cljF9iTw0chXiVZKit6AWDr9bSn7zu1St/cyo/vDd16RCJrhLbT8ls9D
Q4FlzvXMBofoUWLmgu5DsFw+lZwgOoetRPq/WRuitLFDnX9eQucm4xssvDaOivMKMl1gDWVobiCt
HZY5sYDGHS6R5R0D1SJ1IcxJuvOzBeBCIb9PadHF0KcxX5jrcSZZLeNAdLEMIB0dw3AgOKTXrRWt
4GaOvNy2UC65uHlePnJ2BbmZrxbBzGiGbOPlE23CHX+Gkiui6FjzebJAt+W1s5t14QgQotrkQvgF
US3tiL53nUwbsr/WT/fH0iZSCNOVR4up4BSwioYDyBXwA84YD6gMx7WjcYSByF2gQseg2jTU9JdR
rqqjl7EqBi1TnU3cituNsYOzxoSI+wwo5bvJ2xwRulBRox8iHDwygSBVXAcvjHo3JbEdPHkg0RRA
OK009ePm0nbjenMB8+PsVwRzBp2ubjyqfOen/0Qf7/4Vrw4LZDMqopCjYwaoIKtPQ2rjz/JjceIW
5xhLufts1/hmtOV8Jzsr+2Pg41aGT7J3Lqd3Pl+i4dtr4KCnSucRxteqVmZ3Il8p5vB86YZEzLx8
gguK750u/zSK0Fa48EsafwXbSDIjBZ25RP8yN0ABsGHw491lxAa5WD6eUbwE9baFpeacNxziQj42
5kW1mFLahhhcFKtcG2LcIkO6P7JxOtN2AzKG9U6Rf/fuOgK6wBQ45444c0UxioqBzjZO9v/0hGUS
uSrUG1wxk5nzgZKsfImrPetEHyDPb2OX8R49v/4n+n8yZzqX/Nzy93XZrxBaHyWLrYnpEYhbPJ6n
eKwfSMMn/T8wvIlNJUMvUF0kTR8ZyCL68yvEoSAtePSw5ewI4rbmhTHWj46IwR/tJmxORcWmurrZ
9/KsnyBkrNqNdFLFzVa7/F36NBFv3odYasJTNAqyqs+yEvAXDV7H2R/SR+ZGZPo995FBGm/5ztdM
Tx/VA/5oqcDHoR2eDkaM+TKhLGKvcvW9Q9z9yhk+nmzBfCO6w4WITSPM/zPqy6OF/v07s8yQyI/Y
QmRQ6h8I+js0YX+G2KgPjCYJQm3uHwG/pzSQlmZbFfTAqi0Acq5sK8UefVd7Ys1kxfVP6XX/92CS
V4XaC2SEH6IddNCewCICmdG+sNT90m5FrA6FCeujuDYlbzUJbsa2RMSW+20GFAvdMe3Ua/ep5bzu
TwHbPam+AnkBZ5AOOVDY3Qto3rMNSlCUMLT9D9ZHkuypVC0xT/B/PlgkfiwDvDBACQaRjiLx+6IZ
eOI79YSA0lqy/nQ/y5iFM5xh2YN5gISTgE9TJRZJMU36asVIkOVGdNOUDUq7k+ky0LWS3DNK5+Wb
g5N9ZJsqu9EVMHryjLtqorvJwhHXxkVbriyGFMcgzTbok4qgAYpZcPzLJPUxodkX4+KfD6FczxdJ
sSwD2Sn4wAnZR7UiYf4EmObbuvTN6oduLx26pLq1EC8vMWSRnepisrc234gR0SF63XJriBaKpv+K
4CiltUdrO46ta8vk9lFIHCtX62Drj2WHdL2srDL+4maTpv+Re6mOcJet1x9i/Gi8qIvTbLaystvf
j2omAKZca+IO2agQ6ilzIYCUxt/W2VpPkzM5E0SP74gyELIK5TkvPfZYWTLd5tK2LC5325ig3cmv
wyWaG0Is8Q8WbnvWXKcnJYGhwi1X13maxisjY61hX4k6riJLEBC9TzrTp/ZWpXzos8R+So28+yTU
BAJbLleJmr3GN+SUwPFF0aHnpYM7QKSum0uqE/d6teFfmKX1hbgOxyjt8EIdWspvhevf9bcsekI0
DP8x2KNPSMrasGErKB2jlZUBlW1QtlyY9HbMaHVmGfoTW9XkhnrX8kCgtMuYxfDPVylbCyDNaki2
520Sg9MTMHB7v4OXwjzsxt4RRlpgSggzyjFM6/zeLvGUaAfeTmxzs7+Z83bi8BcS/hj2XmFmpkXC
LEDPMdObPz2Zpu71DCbLuXia1Ch1/eKoBOpFJG5keR8UcoS5PN0cjrDICT+8hVvMQLAf/ZbtgWqQ
6UcP9GYU6VBYMqP5Q1zskO17q9fzh7e/2q0PfnBbzB+Y52lj8+4klh5FzX8EJ9NOJLqLX76Y2Wkt
fGX31UDZLQfH3xIGpX07oc5YjK9ipCP6o9zz8Aqxi7r99wvDgXWFGeR7VLg7GjiLE1HVxoPKTiyw
XYC4ILz2E8RY7LCPZw8z89+GTe4TeI4oGakeTV1gAfWv/Kgxm7oEW36cVanp9WBg5wGIuZECvO9L
Yw6fdTBCxDVOG0hb+O2s0i0oJ+hQ33Tsd8NUwsKPbd5uIsfWgEtORyZ61/lGfOrKEXtM12qjF5CW
2l88T6nJSKnHfbAKKeAcQ+AJmH+O/vdjovFqcNThe2/IM1XHW795azytZMm4q60GDMtgBQJISgK8
20EWGPy6I8LtpJxhIgjzSMe1pzfraAgSMF0Pp9XgPI/PpQyim5+iBH411OhOXBSNhaPIcaukKOLF
wvhI20rYgaqrWnrTuKoXOGcI44XxZj+B1ZbQxC986QdE7pEnYDBVAxvL6X7AdUy1TWBhA4tV7JkP
ddVS+/c8Zp9G+eY14JCTrCgeVYu64qVsdzLDI4YHt0o15NYsVbOUq+66YmWy4JXE3vOlVaBQAr9n
jEQmRMBKI2Qvmv6NWPPA+HoWbHvIlyTJiBo7qNbqmnfTfXsNA+LTuKsPx0ESEFeuFZgjCyURfAgS
LFFAQqh+Dt+UEsvCFprUh+jw7+aP/Y3tsffeEyGuvvgSOO94PENH3sQ/7R83CdEu+7gsfu8upLOu
jdyZUNe4AfOwZgrPs4ltWDpkbLgMruouOG6S3itKFiXGxByltTbV5bH+p4qTQN5GDQUtQFJbIYpc
QaWuWPUusA3qax8Ca30J3VQ5RRm4feaWi2YD64A3h4Hh9HTeGCkj624cfC6va+xkBO7OC+KQVFys
sU4rsEjBIeoM1AEHPNhwrcKFAmE9/qfOjfw1z2dEpXwYPcMmjC/55xcoRUr6g3eJqr6gPv3R2M1a
ff3iK2TJkLhbwxGWn/wsy2Fx8VMp82/OhnCpr1JPkyzM68cGIo0a5XEF8QJwqXkuzEHvuoDfGyH1
rFQnWW0I0yG7NThCqQ7wV59i+uMe91Rj0hwURpFtL+oFDMLHldLQYwmOd5ZM6Dm04MPOQCfJTpiv
PXxlk0kqjBZcnGz6YwwZ1SuS54ZaW49v1Tok30caZiTBEtSfW8oX8hDLRYBur/Rx8Eg1/r3II0zR
NicN5c3yFe8+a7kfYEzIlZD2vxOwK1FP2DRJPTNB0LThOzqd9XUA+TXNAhesnlbyyHFqmXXqaqdW
OKMyUh2MDiKXJHo+/Ni0ps7YgTWYKlRkv+7Bq/q6/YZI6m2PTXUvwbz4KFGo1+AizvH88ZkxG/9J
w2CoLeKVYN223rKGFMI5s8WdpMnG/uALyzaQTBiYdK9m9e4YE2Q5yxTAPkKf1caO12b9MdN00xYs
PN1e0ThpTBFcYA/IlncPvboty/T0+S65ZF2yji5/XpG+jT/jzVH35zIo8q7o5luOfiNu5UliZriQ
1yTdREBmO4GSWs7tCA2kJ7XqBTj53d7es2UVf//RBR1YiVO0FJlvSJsI4Z73vpVwpByg3nBsrC3m
IAjhp/IqYrIws5zOztafLeWxJ2pz1PBCYw1REnLX/IZOH5cxpz4xR9i6aKS38LZQ9HGfJjO7pb9l
WlwUQ8tpRFb13QxPnBrEyTQEfyrmz4xyCXtDeu3eHTEZGrCQ9Tw0s8cwMltck7JzPnO/aK840dcY
BoKTZTaxtfa6DmXXvwYLJO6wsXCd1nk0ameL4ZoE77XvCkiyo9+gdxhd89tBo/VX2YyF83hL75dh
84fcduuvB5bAWZcxz9Jl70ECTl3ByGIIg8BpgBJlBQoabMZw07XsX/cOxA5VZIYOqityFggooY+7
C3nQXXR/5g2xZSXSoxd5c88YcGznP85cUBvVgKB2CDGVbPgYkNbvehZhuvS2DkYRS2/57gLHEB7U
p1y5HgAa4+yg43QgQlOVBctmXayMXl0VJvOZScsT3n4dqh1Cir4YI8zyPjPj/rZZ+sdSea9Rkf1q
WWj+PkJiI2VJt0NbzaW5YqcgdiQQWnaUMFGpnEMEMj8OPYF+R0zDozgMVCBau13soubg6+88CLMH
dPSNYnZmeK5hPEsQvr1JWkpzj1PL8e1J8Ye8l+qqW7QEqmSOZ/Y1e30we2f1SwzFDOGN5sqfh5YX
UsQx+rtJB7Ej6i4Qs5o0/+34/x3wIUe/gUAlhfW1Rq1YyCqpXMQvB0y7cHZ6pfM+DgcXdAejRC9l
gpVTeI+4tctFd4ODUNnWidkjxnGV3RJsJppMbGsAB/8bZN96Eg2b050CqHXOK+wDb9TwnF/ZBePD
QzuKuXUxy7K3AEFDRRW4kZ6LjjKD8gIJ/aD9iRAXE9QWYFtB+Qep8IAjVYIf2N34tdjsQZXCEBSz
3F318nNnTF1nrwTLOUc5wnJnhXFbocKw/pi3V6V/gcf4NnGRWhcQE6G74zCmKF79W30sxa05BGm9
LuBHbFBOLt/zitFjk5Y9NWZvAMMyKcnz1XxUbefJkX3K1dEQcc2qkr9iW4hamPXY/+JkzzwmU1ul
5AkO6j8IAqmEWoiN4SuqsJsXXAmj/IvsAZzj0PeNKZukHaiDywofKhhKVjfBj4EEpTV7VjOp49Qm
TfmTNCjNmnXDUTGQUs8xtS0EREYmQnowOD5C9ZFRvFzHNquIODG/rzBAtGoUeGV2Xu6LkVIKcf+O
h16Zvfc0WkTaKr4E/c7UYH9Yzo5ppNlSAfNSDvC697OdBIQK5REUUvojax2gRu/1Dr8/49rE9y6E
5L5e1CTlwDE35bjyRM7Zmf/kDRDK4o+tLVWVxaveX8VzvlGDXqUmGJYT+ZiAAAq+XF0pqGI=
`protect end_protected
