`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mllZavaa3s2kL0m0zDgzmKJijjpZFuFUNchEeUa2gQu4X1LBuYp0QIxZACGVmHRYaHo+cWiQjDKh
hRduN8BySg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ISKjQeEso0gXh1qZgqf5DcnALxlMz2xG2V/1Hu9MD02rxHhFiSsOCsTPL7UEEmMJueDw9Fewa0TC
+OGoF5d1DGfOWOjA6cFNw4oCRipDuwgcczSJNN8RaL2foFCQcn0GGYQuQtn46s16dGx0T+QQoaIf
a0qzVSf3kpV6hhB7eCQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Re0nmQ180f3uadsDKAUnSSJISkEaB2FQmqT8TDgcxfZifsHN4u2IIiANOuYAO6Otli1hP6pvg+Mp
LQW6jAnrj1Dvxb37oStJ8FNQSrGNf1kEyL38mgfAKIq+gPiwZNlkxCeh1Ivej0DjyCdxF3Q59BOB
K045qt9THdFvZuiRp4nMm3pgOyRaLzuetZ5DfcboawTx9dF0yQiR03n3D/u8EeoDKhnEFlQnesN6
Jk3VmXcrMBNtQirc4O7sPbho3p3hZ9cgQnrMQbEoZxj3n3sQ7pNpHW3FB9rDzW8NViO5QPipQHRS
8ni55JprfF5X84OkNrKLA4zzZ03N7meSL+Mhgg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cazd9V46ukKwGa+E/V0Qj5l2dbn8uWWuZu7N/TD+WpiY1w/kN3DhAOKCMofggdqXRNDTQ9YinaLi
IL2RN9F1NSC5UaCWKWSfRagSKg6+mAwQvpMUv+srPANHuxRHnpFuob6j8Oii5UUWjFwvr3gNoGN4
5R9D3RzUfydgetV9FRc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XXTmXdNRj1Oqv4QQLdiLI3Hi2tFkZH0Mogr0z4qs80xX1MorlTEkpMI580Hz3vjOztZwaQq0CprJ
n6icnx+i5+yjhJxdpfXGs68tSDuCu1+VA+slo0GRhBAWNHmIaNPDXecQRVMAVLT93/saYdjaYcg6
MRKBGGNruwDSc+2KyrfndedUemRur45VTvyKmdJoU6ypMfFKOf5QEWPfXlG+N5BUgDVhq/cKOCsZ
CRX6JHgqRe0Om9iPqmOOP5T5FR1HiKwFYWoV0NTC1nP9OnIOpthU9d6p8dYVnj6H3LzSdZMOgGC+
TpLtV82EqVIGHOmL10L/IxRwhlQCfvGUQHbH9Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5808)
`protect data_block
ZysxnBVF1eioPStPAjJ8Q6EqmIMr56RnVoPUwfAFjAMsEL7JREZ4UtEklVmYPTega+zkFeGO0D3O
/ap5ywUyoVn6k6MB7Ran7HUimtlRAg9fXlJUbmN27il+Tdij0IgAfPda1A66A1BjPLuSVDXRzFUz
xozAm2pRbmnDRn6INE+y0gzqHWRtunL8PE2EcZs03iM6abbvKyIuZOVHHm89tgU6bWhxrX+QeqI5
MpklhUTP8QDOsotKTz2+rRZDPHjo2VBwuaM5umtKo8Y62cuLnITHv1kMi/nGyMy9It37MvUbNWM4
HhvvOZXPt8lSint2+abmKE6oJQpIuZBGSI0BUORQnS4RbWcADzT7/W4+lYrOQN27ptupnSKAYVP/
0vTzl+SRkaNNq0L5XS8rtgdlXA+8ejpH2ftMvjlHF5xk+wT0B9QcEx4KMrB216ueBwdwgLvaEQJY
sJMGIfzn6yvsf8XJxS7r8SQnTng4O9uiA8CsgyuIimWF0xo5+AccqR+ywaS/U1g8MSVbTquEg7YR
N7aiaj9JabMWo3U8vYNdwrM1S9eYlTADH7HrFsENl6vq311cDDxveBGbS2uxUY9Fn/KFmkvKALDW
M3Ws8f7fuGKttTSCMzASsll4t/KYmB7NK+cdRAnPyZwyN6alvb8VQuVqhLgap/ByOPG9K8IzPrJu
sI0ahvqvFRo6T18NxPTBtgd1rfs0YH/KKX0ipupgZo/p8CJRfxP8XgGbgRzt0oB1LqNebzi5LE00
xyVB61Ql9Eqaqla8Y1Fhp7qF0QU1y0ObeAQKDDBJua2kJsB0Qah/YmAIUumSH1VtgXDU9pfcDdnB
zPHn4w6fPU5sZq5hJZ2rOBRgjEtkUCd531u51HAQCmjPJwOr9+r2KBX1NzTau2dtW7ZZsE54spZO
tPCHy/C1JYXub4nBP2l64W97bvL36EyJ/JqBqhG6iDauwQUgRkx37u8mIOJP6L24l/5fa0In8K/K
eS1nYlg5X4X9J1tGofbnzb3UIKVA5uc5xvDQpa1i7AU7idnkBtLMTm4DdpWeMxH4u7KtVjJs6yXM
jnc/hEw57Jfko7X9Wf4ZIKQ9RDHcxbcjaVeeeGWWUuf8yaVUwAxkoRW3l1X8PLzHFDOUyZs27T11
RZ+CU+SmGCEUSQDb9uSOqv1d4DoitNEenY/pYFJAyTv2TsmZsme2I5cIVVGG2N0C8IZDQ6Cbpxi1
Xrc2/4XajQ32/hnwpXCmtsJzaVPPAMzR9aRVKjl/Vm0fnZL3nZ33F/JBjNvnsf/ca3QmoDHDzw2x
9mzVpBm6KBIAej7RPKKItclUFmQGA1SDYHI2oowyv2RwGRh1/X/5QMRB3NdrOoHTGboa5hcVONCA
nNhEGVvJqp4y9/biOn9lrOWlvFtvPa3qIzlq72d0To3mXOLh6yPYz3dIqBiEQFx4ZMOUsyhYHhBJ
AOHB3GDOzFchyXaePfRa4FAhL/BssAescs7QaV+mdoOLfBW54dTysmNdpxRFSo9JpiGorxfyS5bk
2/WLjGMx0sShlTeDYrbNioaaLO19Cw3QjvLSTPF5Bi6oCgNh8x04o8niL+LKtcFexpQM9jd7+4vr
HXCYqZbgExeA4FGd1Cc71Io41q3o2EOuVQJH9Lbd9pxXzIwyrg+0UQP7l7o1o93ypEHJbMyek7G8
Y12UVPVIVqJVPN+pm02Tt/lJ47ziqeQowj8FeRVtNNbz8dyp4Lq9Qf45StM4Mj7njj1j7emyloJ2
DnN+jCwJae0v663y1qjNsDtFeQ1SyYnwuIBQww1Sh/cRkm7PSw78Rb0axPv9ZGXMTM/JoAw/ySMV
G5RKu0avy1TsIkxy8Y1Q4hxdM6ldzyQ2g29Tn9MnvIlAtkU/ly7Twn4ro2w6lTg9zy3/5jccczta
ru+C5Kg+w4luADFD2S9aLqSaXcqfwBWYjEOC+n0LllqqjdWTyiMPqfcgs56cOIqadOU6wGxJPcUY
SzHUXBog5yLqgZBo6r31M10DKWcZ1xQY5XoOAQEvBF3jza2WrBNYaP49/YP1phuPIyWXMGfv5bE8
isCj+KPlKcI9KOKp35Zh6fCF8omoz2xzgY1a/npTtbO+eOuxVFzs510koaSEr+c1k1UA8FjdH7fF
KVG5oa+1m5wLEM8YJc/MjYvVpLmaCZ7bLmnkDfGfBpdaDmUCGUmu4gzLqWdHVNDMW6ONfiduwYJK
YAZy5uH+I+TUV426iZUvUtcTFIEG/JkIZJbLrFHzIuAiyoN4IMawEoTMZ3ixjq21ITujDxlkbTvK
qhRbI0jcWD5grrMjtnAsOWHS6Zue6zYjD7EhI7haVb4MAjuvRnGyD9/nCXmVpF7zeRvGMIuJQiZa
lO0oQNPIaOkYCvArGbLREQzzSs2TqxNJjJOvvQ9fzYPhPedVROOA1EH0ZlNKkdrhpXoVH1iDn87/
ayyjOn9AGJHQUOWZfAc58TFgSktLxonUzhxdApCNmD0gdwZNBLGGdyCKSpPeLBFDHKoTH8/SnhlT
MruaiI5zwvsEt//4AbSNGrDvc3bGCfwje31ry1Medp7GcYshCYHj4Mx9xwwThf4CFmMoHc728/93
BQteH2IUt/LNZINE5Gtj0EWeTGVvkkmocx51VwEnV+mf9oENc0TWYtPGzfvITnsMrtdEm9PPeJBs
RYHVzMQEFfDiYrcC0CE45/PqO8YsCWeVRcfGdjbShwPunYbv9WsIey8O79Hvm00Xko1Xug0ArrOc
MYfm9jUSvPUD6GPeAiii48AUhVhyxQecXNYIAb3fYF9jAAgW6zMKVJMpgsrMWQ8NHjQxJo/tLsEA
u8EQA281v0GQc7iHJPGwiFjWquxqnHmuOow89G+Ptv1JFody6Jv7CdI3JapXCLs1NpS1/CSBoB5E
J8ZCCGEDt4J5Zw9+9V+EOAmWxw0skR6fs3aqOpk1vk0QkqcNWmdRP3RvWpIcYmbnhqOW2tOeEUMt
NZxRPCFqgCxd3UBNrm7776A50efHkRt6CZ6DZ5hHrtLuTQMzHNiJUy0bQUz5/jWNH8fY+tXUUpAI
PVdFRYdQaEP2tR8GA+L27moJ4mkispERA6yxx26gKIINjECgBtFRIJ5TLYyHhoBmlA7CCOUz8b6e
tZNFsm4mCDmQB3/SxAsdavYNo69QqTffS8b3NeQHWNSggX6+4euZpN+S8sAkUf7LNG+lh2n0aug5
T4QQTLNNQUTabJRSB/h8mEPgCsBBSuDBPlcYZXzcqxf1aUIeB7Rrv+je1FgTr+ISvSlgKqVRg3Uk
/EGTYBYTPKO9lKX9yjp3a7oBJ6JPi/eJ5YRHleSu4pYG5oGgeOM696t1hP9Li1sZ/Cm4DB02PZ6k
OvzZTPO4nsMXfnSy0ZmH6Lr/fR0HWdMdSLskd2TiqAdLTe5e9yqiOYVCSFV9XI8k9p3Xzt8BIZtF
BHItw7DHE06jlp9G+Jc/3yfUzplSuYrqaGrq5T1WP4wr72oRJB6UNFr2wzFfn+NWM7gp+m2v2jRd
N6VC21zlDDuN5MM/HTN8YelSOH9a5uoiA96j0LlIOXYewE26xWEXn6VuRgdzCd/Qv8gKrNbQMPMQ
JCtYoTJUq8WRsFejPhTexqS8eHM9/hD1rYjSAPYwhTcWRWzc9PWDLVF2kwV+zshvjTBqAnWb+Mbn
+yq4ryymPkmPQI43z2r4SYVzT3Eip9rzxph90DfmB+Qah1NMAXTylbVm8zlkW2olt7ouDLRC0fB4
3oDNqY76tS2A2VkKort/LY33PNmtqYlqbZMnDoMSANYbfMmLMs87YJJQIBnbmqkEe+0YNNtFKCUR
1+tHIyS+B5+DZfD96XOjlb9cM55O5jeaFy/40QPvuBDTF+oxRLFUYdTJFFu9DN02636bvO5cRxib
itjI8LXHdERpi/B0P7PPJBJkXpmp6kwb1WvZgfYWU4mvGketEAm9B8jKRe51y9030e/f9KeObi9c
RlmqdkiaGNcuLFh7wCSihC+DR60oNSNPKt2Itdbk7Ixi4Gs5vw7upAn0/itALtmubw3JQMMEjjbn
tafjKQ3q6ICrDy2m9GeTnxltLVPbsFfCQlrA+mXmZCDd1T75Gmnxa9xUzuEZzVDdwrnxTJEwzpEp
Kt8AnMY8bmLolP4+VdE8Z4VAkuZrn1/6I4nUcjb+iaakmM5NiOy4Q4nwshoFlwQWG5mPjYFWKIuU
2tpcqdhXsIpeLJifuqjR+AUGspPpvV3U41gY8DlSHAsTFszxUcqxJZvM66DTKflqqwmEBHDugyUF
bjGpdlSM5N+yqJq+l/ibj6+1s5VyUIssoXDwE4pd8IAVPKlui8xq+KmymefpynhrLRkXoi0WtMgx
UCM+cRE2kRERbpGEIQ/lvXDkWAZ1KrwKpkf9tj+wGPwSOmV0+D6SMJiUz7HApFvKAPtyqnUv2dH7
/XqPvn1BSgER7jk0J1g9EwTbAW8d4VcWVaZfRNj+pSlUuYlYC1NNzaWnsOnHdOb9/yTHd7MwjsHV
ukhb4Jbp7YAC5CVNZOrBBwMSQ6S717kUHmthYriHdOPSsWNjc3NE9viVbGtkVgnJ4XB5cZD5LKiM
Vrt1M9iVJaN7AQcEm7TPgvfnqdjlSwpqj0NGYtnH6q63Qkjq0+XExmg820kwd2Kh3rXChlLUZFvw
83oIwGOFU0UGAsY2boSA4V5nKp50qNo0dmz1HYunTKc4buedA8BzMCEOjXFXiu1lP8NBcjxj8Dlw
wJhsI6ejbCx4KLewHE3hdv7e0Glz2B9z73UvqBhKMMFhvFhGiD6bfBZyZMb1E7wD41Pbr/F8uxzV
ED32/wowbvJFpZU4uFJOb2QcgZ2ZtQXsEGMoY7FNJ1Q42qbulY2b/NqErKqscmmd65aUTGPMRNnS
5sQQwJ3IqTnsIbiCG+E6vZ0RHz3ey/DJuUUYz2wzpnSCapz6GD4h9sETvhskqAUAAznGU5cdjkGp
m44vwM5WOk3kap+oUwClWC+Tmr95nEKdwTZ3gYEOmKlnYBhHljmyUigAbif/8FA6UPZ1U+gOWNNj
LJIQae7Qniidhrb7lI7qd+7GHySqteZv2dhZqsWCGF99ukp0EjY8naY8mqvfpDM9PaWOBbKMvH3u
FBlRWvh1Nnl4r/QKexeHvkuXTh+urPHtIH7WJb+oxwqSeB5jv/Q9Ix2MGZPwfK9BKK6Q1Iifd58q
/X+6XTYWQK2UgPlvShdne0g/2HoJIs20WNGlLWASR+0vz4C+YoNVyZufeNqaXmtXWsoDhvdgPg8Y
USLEmcavIJUMK/DSdQ3hYnlyEnTuv9TOTLPxdY8P5FjUj6MvO5Dc4KyvbJH8ElZ2jbe7kczC0+x4
Zssi6agTFVTgj2ZEgQuq4yG+b4yDN2FNYf/YDVbb12HbOswgj7uZVCpibYBlbv0/A6I5dvw8/2hS
VBOanaHjdYS4Yrci2by2YNQIOIQJPgX4Y/v+epOs3YH17JYiX+EdcNWYgWwkQVijwTzy7OyfrT9v
EnnBUlCdDvhSSc1eI0mY0QfYYv64TxH1DH7Hnwu3lBdGTP2cbpk27lmaif3ichGuInzzlD/jqtTD
IDPVvVhTDC+0thjYcGGakoowsK1HpDJLdbSHlF+wJ+chcF491ONszlWnz3JIdm5bBnmtVox6d95X
Zul7taoG4Gkq2Z8JxA8jjFPicMVO4uM5yXRzjjH6Y6Y3HvFdPbmWP0QuT3wy/CM0lTRPTLD23XcX
KITX6Yjdurle08WK5WZz3FOd5Mn64j4IcpjOJQOoL2mHb7IbU2nfgHAdcbBhB9UnoTGjHxi6qPG6
/25m5C3jovwlV+3ajeNCoKKLWQn0ziecj3vwWWu0kVSug6tXnE7VVBcP444LRHP5GrhTzJqkjEc5
TRSqL1D8qrsoJS0yOV3Pvk/UpQE2pYJdAnzFrRaYnxpdJ3hh0Qq+h/OGru+ST1n+8GK4qtqdid5C
VQA8BCaqNt1VB473OH46Bri6q+nIidm58SNVuEQkUQKYtoTAybbgQp4w50fCYuzo9uzGygDlA0Ax
33Ol6tBpBL+jSZ87rdj2vl3woNIc5ls74xJDgyuJv00L7sI+EGGVMs9PdZLpoGI4PE06x0MJcGxC
JzhxLa5x2rFfEsCWFXbBSTWecV3dGQO+xUfN7ngH5pdYbkbbWZy2xg5MfanfvKm1kpO+H1Rke4/r
owCaDBMRbtE9LmX8+/dZu0EGmOToDrNLKKySzxaQqv+3I60cKl3MsDB9d9GPIZVS3hdja9nM8TZC
oiUIFakJ5HrOn/sk4h1BJ1KV3y9IcrdGX7dPqkiHOpMeOhni1DIqJ0zSLY/qj0pTcR676F8fYIxb
WZYpwdjzzFwDxHBLScx7cbDf+HG5jSGeuD5qrPtepkGv3RZgDZMFC2Q7ts4ifDUYJEcs3Bz5Kwh/
3N1KKCSBgmNpsEuG1RG7oJ68y0w+GmVntNMsPCDZXwMaiIIHa+N1AiicmBv/9bt4rqdbKfQeg7Xq
8NOo5taan+lZxyZB7VvgMAZkQBpW7YTJfrbS+tOm7Q53OaEAMHz9EU3xdsg+fZWQGbZd/VwYBt00
fxT2xl7mDzIxj5mmdNuYZwrj5mxHFxFH+xI16WvPHSLn77MgQUiCHp41zzB0KdqGJEfq+a5M2D6y
h2jhbgFOKd0cFKy+gAHvNMf4455PK/kITl43+tGkhJ9KZvAH7JDBzc/iaSSg+JiVXjMNOnPL0jT8
eorz/9bh4/ZUdR7nuB5e6pfCWq4jRankE+H9ghQFRnmOOt3wTU5gWognrRAb3FFOUu99jteMSjs6
0mcYsf4sYfjqhyNxvPLcU3nBruvcUxT0kW6a7RQT5vXVIJhU3iVK9HHIaLe+lVB2XOpRKfdsn05E
XJpv1ppH1tYwSrBvGaa/Dvq4ddS6sZzZqK9Is4oaviv8U2UWaqoDSrNMC5rb11RKoQ3vUdT0LDga
QxS7pj/YwDTplT7kGtsXlKP+xbboeLZqJOLTxbud5xQ9olu/PEcwbSZekflS+jBcHZLFRMDA48f7
UFZhHJjToFIgDnm/Qjq1Ewmh/fyXbMfoBhKe2U6ncPCIpDU0ksqH9y7nWSxmdSkY6AG98GV51WgY
LiT0n3jvKqVK+sSGUnHszyNqRJcY0JMncLwUoVs870bVSjkfnWJh6a77Uez+duwS8AIqcVGwp2RI
xGK1gn+YJxm6E81fIp76tKewVYQFmC0sKnmhQF+n0NKiklACnB7u0eOMZVoWK7a+T0zAfaNtZDqx
H+qaWX2hGKBqQVUXQbnd4nxnO3v984NLtBhxnjQwxGY7+4iy1CHdL3paO3zH4df8GxMBZIfD2zv3
VOihihzXuUpj2hd+9Lhifpu2nVv3/M4+cBp82o6Gitt6WBLId2gB5Qf3b1aK8hfn9/wX5weHUOvg
gxw9tbIrnUAT+9QzVeSwwIbK1/xsuqJ+Stnxkw8wdreAm5jSOI3WZavMkc0ahDBQTW4qfvLwr2d3
qcnc5GQLUurgpBjZUlRj+RWZy0gtc3968sC/X10YONdXvpLkcq4hsGUFjcSrwcHiop07J3I3qzty
zlyx2Dz3ZCcnb+birMCVzK3QuYg4alTDTvzbT2VhS3FiPFOSRCTn7kKaF7TFgwwB2TxnbckQQ+nl
2wwcoapGM9Bca/9zPd8lcSdZZy308nVH9mtT3lp2eI6V5mMliRzcTvOYyT1fkbQmnYoqd8wZR8eg
0dAurhF//J02gmxJPf0/MK//OsYM5N7vxpbLHOAhTxlRmPJtLHtHYPLM2kkxkAIHc1b4
`protect end_protected
