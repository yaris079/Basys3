`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BrVkrGATcP40JMjnflFSzsUkDLJxCQKwYII/04LtaJDu/g4LHhUJsRCZmJqAO6/o5gywtv/s9gcR
ta0+wLcpfw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YkZ79lFhh/sbP2V+Ebq7oHD23BK4FZmn8IBNmdzboumPepo5LjZ+KI2JnZX8nDAwOziQ+A+S/De7
PKSTgILU8DFMpQ0UuqBrKIDRfJx9RrVBYrnlktSJIarpVk52fBVj+tSRycuKw5dPMzQZcPz4bTes
7uqjRBAE2JOZQqUKS/k=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fEjBIINF61tiW78QduXGMA7sCugkYG+7MnRG1ona8L1LdsEEgBzo0zfh5xKHImSRIsZap6FI7VZA
SpXfw7IE4d+ASRlWLvvAn1yyeDcsXZT4b0u4jv+RbM0mUFrOPGhkD86X5lwhnqHejFWV5L1LpEcr
3y/1pA7+0X6Tz/Oc5zzM1mYgfAOTpJ/1itkC9STFZDvIuC1K0IacMHOkSa24pwtdFChMDXFArA0O
hVPHH6JKrfp+UyqQWrWBRBxUGLDWrGQGOTcl36d6f7fjT7H1j/YerHEwFOjBPwnzUuMsDu2390Et
Jyi1EkMCGEk/+OwQNtALvaiGVysdqUzJ+f93Fw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jX3OFjXXr4caqb+nWE3mYv/r+paqgg5xQucoA5+iQh1gLcaefPG+eM7bl8QrXYOXhVK3RyaG7nuX
X1z8S9N+gOhmtcEcXlyeRByKj2GsbEZTFkhr+iiqXbzGw+akq1B7HhU49i48qKvUZVPpBwU4uKlT
2PhuT90lcN35StGywJE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FqZ37+mnTUmjH3ATPN9/rnfT4Znh1mF16VuE0ttlXlgPqx7AUHfOtubqQPRUXxtiEiPlqe4RwbR5
1tBOVkl4BLJclDyFsvLsTw2tFxXm/rncVnjS0YssOPIBtsjClYEDnzJu8Fck7lJy7BQft9on4vMv
rmAry5zpS/o0L4bus5xHSdLT7ifdGyukdISU0J9cUoa33BlVB+HSGDFi4oYmrITgKVzyN6WUM5wH
t0m7MtdxQ8f3ZKMxHCzQXsflVbdWbDWw4Rm2yL8E6tw5lWtMQ878cq1EqXVR7ERHSd1xPIP2BOOW
ZaD4noHUjj8dTVWWdmPQ+1EUAR9vi8y7PZ2dmQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13824)
`protect data_block
rhDcijk/KkajNtgwun+8AT2wOErg2mWcEdk2Le7EEtvEka7vckhXwghS8Sd6XvpVOtI/4z4xw8gG
6f/svbNuCuIYYj+s21VRB6G3j1UmIDUeq27v9uMl4CRGtgpLu7jPzmKSbXVISedsi53ubhxB7yeL
WBSoYwk9EvUAix/ZuncwlfljmZ6/IputBGxeY4LzygVMpZZ6PRL3x3AWg3YUUzt1E6A4miolKicZ
YbNVtpRdBUGxv/lPpoNX78HQh6A/GTMonifB8ViTezYa9FmWpfFnMpWDlhbTWu5yG9NXoZIOvTbP
6jOMMKRIH3EFWT9FZeBggEUKvoyB+FXEtn/QZTEC5T8nlnRpbmGbPknm14oGLaCVqw3S/ZxxdOFu
Y1plmmaooCJhknrOtWEXhjIcaFJFsbmtQjryuu+gVrAXuNWQ+3ISCv8y4H32nXXEmknIeO3HU33G
ffJT2PsEFVa0irSMfMdzwPV/8yODNj1B2SU4e2W1GfZcZQJiueT8TUxrnApeVGaBEgnbJuAKcHUh
iF4OSGDCIyQ6ibRFqYe9ixYoU3bbckQRiL2Db3v+6HqQroLzMIlS4Lp2abeRusRA49uHtQRmJsBp
3VIOkZe9LqTuY69ebV8BhH5eJ/lWRraZiCUncaREIZ/Y9Z1hceAfvcX/8ovhR4XVLLNd3JmMxs64
l6Yr+4x9JEhRqE3kxRpZeBMPGRjXOWKRvxW7v4uZ3YI6dmc5GthGBrKqgz2rqu4apxLIltcEcPXv
7ZLH7idK3H5fAE10mnbVBQ9LOoOvyZ0Mkz5lE5F5llD7/oTy0+tNbrLCa3l+KqayzGZFnNh4i+zj
nI5Bf6SKc7yxTKcKtnqWMj6HtlV12uuQ9+rtnjgg0tHcmKVmqrybpAvtuwdabIKwfChK8a7U6v5m
PE344hjSLRvznQ+GvVcV2hvQFFUITWkxRQFcyOQLMlWXVTQ864PXVlRot2lAe84pkEsJflbzUv+6
+j9cZq+c/HzvzUR9DwwHUf4DLAWLUpxOJPdaoi7N6tfNGjPTihW0UrP0+zuIVMtib3y8kDMJazbd
V+uRi/gkJviZ1TIONbiAInUyj6IkOvd11oZ0dl7aFu00AZ9uR+MCaL2gIUGIMQ35c43jgKI1Lbgl
GXc76kANKGoQkBkQj+BxdzKWZ97+df6DcrZl5hO2UB8+pgAG8/vqg+WumBJTbuePEIPUhlQLNs5S
sNCCSbmdewT4uV8qyel4+DvhR0ZxYkAN2wzil1tMnci5SRo16Ig/x5NB3CAPe21BgPSggkYK0GAb
jepLY/1jfvAQpw1GG//Wo6A0ZopgWqMpkZBXP2VNIBXynGYFPWf91mhnKdGz/XswDA+onlRcC/SS
qjppfXs2TrdimUu3Wst447e/cy3c0/cunx1raHIrlj4pgqhFmhlfEA927Df462e57f6HrTrf9NW3
ENawuTC7F1xIhF7EMlo8qZ0b8b8qItqOEMfEUaOY/b0OgrDIwD1gs0lHtZfLU/wtTXhW9SnQZL7V
HLyT12a5Ql9xqi3l4VlVwIQBeIUlFK2dv7th6kjB8FXejCDxASVnkK2YQo8Qev87WQjemmH+pCX5
MFgvwzKL+0k8wazfkuzb08VVGMHUq2nUHLcbLXCJOnzV2TXCaOV4j2I/5w6kSjhARtffrmlhpwz0
BKEDjxYs4FWnYgyZBpTge3f5S8rknx9P4up47wurHAjvbD0GwH6LORPa/4DjNmypvLHqXtjZjffu
XyWi+3rco549Wtbht34MD1H7JCAHqUfL/CffUYApGfikQraUeW6NiC9SyHoE0eYOFKexXXB+kMFn
oCDYXGnxvNqddmAIqmzsuMLdGm8E516xgCAvdcq0lrA+cwHCpEgH24baGgzXsyPfNi8vPMOuQ4MJ
150cldLLcqzg6yWL8JrIUbByOR1nhHBI0+FFu5cO85kRLAUStmDxYXtOy2wHmYiOkdfNlMGKQmoD
AYQmxuXy6ETPJl6/tWbde6uPAhCYIPksNM7eJmE4774Z+gnRsOLvhva6S/EADCH+kP3fjurjqZ/h
kWeNCl/69DMH6xxTiCNHp8aPpHLP8G3jQhjP6wpPDp1beNED9tyPmbedzd72eZC3dfUKNH+LVhrQ
PTtO3gy/18epgViICiK82fd8VHTxEmcy2Z9ejIbB4MhFXqd5JrjHGm4ydFH1QiuvC5ko5/A9Ihrb
G6ViW+GHK0jgVlWmYGV/JbL4XqJNW+CwgIVENy8yXvLjDcKeXR0b7SplbtA9kHzb9hyv6a3oUMQ7
MGKB11ek+VYrljfb4HT1olpae4Q7wtwKeMrOdQX15dGGRxZ+3OS64iAevaieUS0+vv65K6/ZJJY6
Ez+KAQ6d59qSzjl7zAJzd+7IO0izLFpK6FXkQmXjnMURebF4cLTovhm12pLIbZ94r1/ql4sS92uM
mODs0X8wlZBTk67/waIiSCtg+hFykgthLBGdltHlLYGQq6002HLgEfdLWDulREqCk5bWJpPFnyZ6
YEiV96kgnAe0AxOOYy1+9K9oaSAVCew6D+jeBomyU2jPQAPUlle+TAStwMpoejRXbZ6os2uKqikv
Axz0OOUbdqClQNQlJjyvy9wdwHkT7Z5Qt3rLhOUEHXkdfhN7MLPk2cfHU0TFeKSENYGVbQEpE3js
y7s24sjBxmP7YUO2eZNFj17IYxfjVGeDc0gdL6B+RVkDIww/KHN8IFamW/YeLGCMWEwgOuYFmWUr
F0bUJiOkzrVJRenS89qMRV5zQ3U7/FTqwSmjo6vUbkm+Jc7gLFg2s0N8tv8ChuXZ3GTuEbwjTxUT
RTYq1IQbxL71ux4Ij3o9nJrCvf2xQ/nBgU/Ao1F1TWCQ+aiTp1s6WBT4oPKF9OToKfUN9wvpP5ce
OCeKzGEiHtBH6PEzpUIJ3E83+Dqja+RS1oByA/2Ew/SmyhKuLYEt6TsV+BqJUa3AGHcyaJNMtSl9
LuDKaCPSf5uT9O4CiBKWPFoKQBgCDGZ8K4UyforPJpODFw+Bp0GHD1Drju6nlzrNg5dU9P1Jh/06
eyHW41FhLh6NFSvRNQVBp0P334MV0AHnv1Y5lIjk7O2wsm9TEmBUXB1ovvoEwCXOGwCcUMGfWGQe
IQuWnmCcMgeK3cx0YQ3rJ3Jsqu5uvJYgdl6YVk74erMb9FKwnmOU0Tj8OJELbM8a7tp+OviGVpWc
0u3EDuZwpEczY44O1yo36avXXaYXNuzZxQKdPKOJiUUVLIRN5KX9fy81VssnSGe2EpH1R90xR3i1
Zwv4cUasceLQmmXKzd00mAHecrV0/YQsvO+96zJZ8umxm9MUkySSDcS+hX7GTDKGHfGPzXJja80t
zufnT2aQNePMRDqMjRrLK0M0XTnkmDZ/hmHfhghcQrDVCg1kQtfflQK9Yz+xREidWdJPaJr0vydk
fIeje0DexCp629vF2fMMmJqbOUjmp7paeO13lNzM9ff4VaDWHJ/u47FI29vU0bp1f12kPNfUIMOn
EQWXhfPgjmFvopUiimosh0KDviLlrmrJbVNCywngBccOuA/MQABligsb/jwcbX3o6IyREr4MQRL1
AGP1qwNxlWKRyRjxfE5rblnlxffuNfzioGHkg4GwXWeHHzVlKhf/4cZngNipeuXfInvAi0DbA2kZ
3YaB/7C0f6FTecFxN1u/MjkMKOlDGoupeXQGW5WSUm6OFQUy73I3xfad5aceBzJHY43I+qK5iHMn
J00NnXsS+3emORt22MqR50jlrz/KNIPHtnAGtLpxqEMatzVbW7CV7dapJqLJfwiMkZ5AmnO+24US
kXhJ+Xolb1O+ksJSIoh/xB/yc1X3ot9w7KoSkHez5HDj9gvfYtdWlLNUzGUJ7BUCK+IsAWnxrJvH
am+EUCXwhvFV5asnuFb10EJFh9XY99EsiW79BYM069ZpEh+2ILAnaZpoYza0QoVcsptc4XFL5Q2M
idoPtoG+jE6it5wY1da9/sLhUeF2MIFuiGhOXEKIlLFvc/3SBM823yxxwtPk3YP83RPFTY9zBcCO
FAm2ZpJEHC7qFdCrwm1a7jKzaNs+6xXoz173Cgn9IRqOqsJEDQ5gHj8ZjaFwgQaKg2gJpvyHldGc
YC/QDEuM9hmJ7aPG8MVF50dPx8CcHKch5JA/nRqQ3sEi/7v7WYF6TbqDHH2Fm+0jmmEipg4TpdkI
MHHpflr68+R5r5ThTPap7RaF6SMLeDFQxgjBFvXvOWMehFFkUCF32ouzuZdkD0eorVR98B7n7V+I
X3Nwbfk8GWhtxWIscLXwtMYpu+10PS784f95TfebGeMT7GlAbjyLZnxVfk+TwT/NZwhZXdNFT0xr
7yMjKPc7HpS+iapZffSe2SgvKdwPURBVoqqw8WCEjZ34UuTB5SKmob+1ZCGFcCuOAyyoKbOv5biW
SyNOC9Fy+Ni+aOwT4XUtjiJGud95RPlOR0l6gSGTWieVLRkk0LwElxvFJr6L8ZDN7l79YyRtD6+4
H7ZXUOo/nCdIDTFlvHy3u0s2bWeTqS/fMrsXEwg9nTsCpVwMGXCJbzCmuBPEbQWQITFzqYG8sFn4
XScswK0WL8/bae0yyHw4LkVjnreEjAl+x/P5vYyvi9fAC/NZhkR3E7BbpHjrO3FcRtLzVuf/CmvR
DLI1ExEtZSFtmXRvqHqixxkGEoZk+waiUcpEaYN08Fy2nTsvbV23xnmsFat+9VUL3YB9QgHRU+Vj
Fom8XEqZF0JIz4EkFL52DXOYSecdxSi8A3GIidRh3pbMF0gj/T/btWTqsEGK09lV2pUMFWtTEh0M
Brs7gWBxHauVRA6S3PW1fvgMA1edBAX2UIZUo0jmss3gf15xE38nLAKJz/VyFZrl9iNGuHwXE9ct
JKmP88ChcqDPp1fq5Z5Sy7VYg+ERTNWQmP43sg5chDmtRs0Uz1b1XIhOVeJjY5IUarMn7jtO9j2U
ikllrIdmvcVJRQ7G4QZ37/AWy8PR2uYYjg4w0A1fZ9QuyjURtl05q4Jl/PoNjnYrA/3oXKgAF26A
/tVGhYS1h6HlITNmPLS+18SecHy71UfVilhNBYs0DpwVUJ69lxy7sPOMAu4nnLCNZrFLY4jw9cI+
zd5KgPyGSI5MPt+qAIRlZ4DiSIpZ8ikxOYBtA02IcZRaJETKuoNpcJc/vRVZ6WyMKmv7jCZvOajB
RGJ5gQG08kTNDTpN9ht36V4n/qyFEspAM8sPsuUJe9zwSiqXKj9mHRXSPrR9nqPtM3d1885lky0u
Gw7WLNMX4zSlsy9O94+oWXZ0tHcnPtSFc7O88olOMCvatkMpcvY7mi91o2ZcoaafzSKgPkSYo0Y7
UzBYaQRIIi3IM+Z8lM1bGMo4NIZVvzqEoyClqlaReryJURuLQ5d1d7tnVhFAy7NUxoVJw8pS0euE
lURxcuozIAiMla46RAmpPVE1/C6QLtG0TFsFBknbha06NoGhcZiB+FWKkzmwx42LTFUoRlWTNSco
u6Q+6vTXAA9dRRTsVaPng1pEkmjTd2P+nLoE/U80zBUzvbq64fGoCrh0kZlbAEhYS2OMwXEp2o6p
A7zRfctKf9dXtn4BgsXqZBvtudNBc2ESeJGfzMALiDVx4Rq5oyxzkinO47eFhLMhObOvlHekHR6A
KmckX70qkeAdYjQfEzUUD42ayOQchd6dMm4V6nz2ju3vq0JBXzCcF0QjBSTEbFEpH4eo+ujG/VfO
3504YCe7hShr0PuoSySqLnEuhNN3LLClFlv/JhUDvLxOcChnqX5v9Vkq4tycIrzMLv5Wf/zu+4JP
+9cg7BYPd89ODLSb5fSyS+kI3bUK5qbeK+ZBP1vj0tqMhr1yBLhnN9iOA+q3xss1+Tt0fXeKbEmt
p5ltxeo61K4MMebEaxhmlC5uVy9jvZumoBKS3ST4oknv1bgyC2+RJoImEuSTW7Su4upYbxYgEaE0
opUNtoW6+ZsMe6vwYfh5wls/8I48gnHqGuYPX/o1A/yCVFlAMQI/qPpNYC/+j+fK4WjDuwRFeXnk
3nxdfXinfXMjko/fssWjj9raMh87qf6Bfs/BtSgGX4JwzFvIHi8OVy+R8MTJwOQR/jEMgANsmtZr
NEAyoXwW01w/8Pac/5xYzOUx+WwFgfuyevJsvBBt/HK3kiR1LHd5H5KDuCbfZ0Ptj23JVHxCkwW4
Kyf/+fs9QdGUIbvfZ0o7i0mTzCA+aiUDXDq8M+yylgldIFxX9Gc/RQkHF69e9/mz9F+CGWx59BWa
OqGNnW61wv2t5oZGljI+M+WczjN+Cik2vJf5N1UzqWO3r0IXtvN0ofz0HbG8MrwrA9spwC90zQi1
PX3bBQ1kthOTb15kcn/XT2AeZcKrJ3RSKQGlBjJ5lkHKEJ5G/07th3j159/cW175eb9Bl8dM/8sK
AjjeSXY8iWT9M4LvLI9hVg8ChnKST5tUHMJexl+auCzqqqmo2uT0/RfvMklTIc4Pw9x+8JA8Fhc7
xIsJSKpljLgL8otwBTGQqy/qPRRN95GMHABwidECWj0NCDzQmUkFuxKFBoPd63fz5R2YlN/+X+lx
fwHp+5duFgfAcSOJyMZYcumoxDwKygNX2o70u6kbPfILS04Z85KFi1BJn7+j05/eH4Vw98db9Vqt
bSrJO7V1BfhYcMlkzEokh/cWZ3ZO4sJmX822yk0nmPy+VAV0AcTWzivgt2j2wOsd5odngGSx7oVx
K5GHlC0+2pH/ghUaN4vG6WjsZZZv0Dhad1/RwHyOV3DMu+3eUdwjRtmjIp+oBTiyNAzFUYhzvtup
M4piWaMTSOzV2n4XaOHupCrMxHVlHhMQTFG4Cbu5zGvL9c2rsQ7R7E1QcMDPNnMOccG/sUB25n19
J4c2hgkCqztK3rtTo84WIcnXXzkYZ6OiE757LaqgKUOscRoAFP1HHf44c22b6CPDxdRhmVPph8ha
KXyYwvcQJFjBIYD4ro5MNivi38i/rtio/9Z+JKvoSCVjpbkvJpWcq0MPRr8VxH9n4kBgQ5Glr1Wy
rPWdl5PHs828C+WS5m9V65nm7EiIudpMuMAoUkQfukUdtvPXCkUVIrpa5aaZkk7oMUnGawdaQzf+
YRsS3D/ZOImXOxPSmf7uJvueKOGsNwptGrFWEn8nz7G7BqWNrI4gonkMVcBq0263yxNqjgyml7Ik
clwhiHVje0S7bVZ0UQUMxPBt5zmvTXQQDsLe7r+YImUeSHqjqFLKn5kNOFqfhU9sl7kON9uC4TBb
FniKGE+fRon/ap9qBP0l2vf+fNFKtvWtXCPPMnY7I1Luc+CwV/8yWaIWZCN2U7+jkOLS72AJnClz
zrixouArw9vaTxF+mbUL4f35YUc9NEnT/F+vD6qJBrnz4kxVX15pS+0Vj6dt4BcVNNgF+9KS+0vH
D2FcK+ip44i4CqpG39rFjgi5l4SY7qBIwigbCbickXtfjnZ0AwiO1v8skbBczq55n0cVAJF5M7gu
AS4TF8Gl3Lh/QhNLBvSG4dx462Q1hvebYLv5giX9yJCYI+AFymNewVg3YggR+oigjjh6sQ91637h
0paSPG6Dzp2mu515lXG8xlmLRKITXOhq8AYe0sfw049fRkOA2L4qjJgGxGZfwFLhJ7wJFsQxsjup
yuWqGfkzB/uzOujxOxBlysh9Z0qiRT0HswCJLP4C8rdN/lLOjfsO+r8DLSKMgpPmym3Qxnq99ag3
cLKgSDSxd33Z1TwfHdPXUGDLWtWyMaCrXy+XXqDQLVrppnsrYU4T2d2ETLp0FF0KRvme9+Hz5MTJ
8pNbWTcEnd+PF2JmhKHOMENoJG0aDhmiR6SUV8IMvRZ3/BNZ+sNAnAIiLl3EMs6TnhQxkD5gdRF7
Ut8a78SkMclFNb4XYfwpT1WRDOESAAdJTXGLGvpFbOIrkXtFHSsFOpr5ioQQf7F1+774VNmqMML5
bowGtrdY5BOiGkh22kTz28+Xw7G//mFiiPJj06EeQwZQdjJg+GNqj22VD7/kvDsABY3SDtsnCVuU
2vNmc96KK9X1FwfFr2Ii9v9Y1JlnxQfbu1MBC8rruE1yPjgrsn0/V7Zfe9M+0kCuw/ungYfu5omC
Ie9J1Dy2PxoFEZxTcBTeLXOvLTKVpbH7gmf6670dJ60dz/3GZHljtq8siwOjKO7orbp0iTp5zfI6
F1l/xAFYwgkHgXlvejfk4INX6KtzPQQ7i66XhZXGgJ5GuVZzKzHeLxLUl0puS/xvnfWN/XCFsMCK
kvKBWT1x2oo7pAkfJLuLSEbUjg/J3YSj354a5s9GGRSswIy/I9cwmTZjndMJIT1yWV9CumlPf5t+
sUfR2RUNOTKIbzUnfGXF04ZZZ26I3SHbZpnloufBkRXNbctcPczqFkC8+00z0ZLseHVtBH2YWV+f
UYrU8gAskAIW274zz3RsW+Ddr0PCvTwx+Jkpy5nkLYHNkAiaXJMHfGGACrXG2Yc5n5GMpMQZOnZz
lRZgRCt36btQkst3C9UCapgLUX0khwG6IjLCe8tPI4i0Hs2cPp827YbJ3dofJpNmohkx4n9aDLRa
CCTyTamN7n+W14v+gjHQLtrD7GBRiSBcbBJ0AjK3yyTVqlEf8FfO6gbs1IWC67dmNgNAXnsZFk4q
bT1Gj4bfpLP9o/CH5F2u4UBvTGaYqi3mVIQjT3mu+hLQcG13LGWnk1TeeeM2AqEkKAWicctgjSPN
WQYS/3TtlQUtn/3WSzQg7FpfojDhNWbZzTXiDZRnve61l2NELBwnz3SVeKy7kp78358/O+kNq64W
fD3ay5qwKnuaSwXbxKZDi9ZwVS6GiUkBVlsvdR9kvggMtRbX6vqz2ARXHCiY47W8P0ElF1OfDXam
Cs+Cy6/35X1lOgkrlsORbLMgqCmAkOfSLSpDVYXrANixd/FTF1RzlYMrZEtGYfFnsAEE1tFaDOXV
ckQOPShAf9uoSzTH0dYhCrenTlhnW9Ur2AefBlg9/2MjPdtvRodZGEPSyV/mjbpPghkuSkfFEJkl
x3Rphgwi+8V7ZnLvz+ceuw4TYjF1p/RPxCc/uSoE6lyPhl8Gswm09dBKQX1wne+MhEyxPOXgjGoO
IBoEXkXqEESYOCO0LoUUMyKSis9XSD9PGhZoj3Md0P7XLERkBoWpltnG+/mi7JXEOJ0OmbBn+Z4j
odLzq4feD/Zo+xkWvzrJoRHuKIY+Ftd8WRk4xxxmr4o6r00+7LC2xhIUKa61+aax6xBEZSdNB1bN
d9GohiCM31H6qscsMoQXhFgDpScinL4ZOq26YcYvIl1jKjM+ulQ0vhqWRG0fYs9FaoYu1ZTOlXjr
qcUZKgw0jGOozU4NXmFYfDWm+NTqmw4Ymh4JA2K/56xjg1THQR4/1+u0Cz5yo8Zu8ARBOxK/AP/4
vJgyou4BW7CwxGX+4BpXgEwjHDRSoaL4B2I0xDymKcnDbPABlHgFvTs9crho/yp+wogF2NmERzMx
etZpQ1ytTH7mY1HkoZRg1hMfALr+SivEzrUzW7PDWZ+zeVflCu5rcvYiv7iZ8RaNwEdeLFecbWwr
qx84S/CvZISvW30wnrUSAbQOmOw7N1sm1OiYX2tEW014s1hQcf9eP1KYgOgujIkrjeHAcsqDW0Cf
ReAkMQZiJVLoibDW7uYh5Meknjpw23frlP0yQpMEgHLJLNHH5Ql6NN7tlxY9DWataXgneBD+mNp7
7jKY4JOweNcnWyoiAY4ceaMMs299c/kUYZaUYdApY0AN7XvNwChrwqxIYuvDkjeI0hFPazjVAcZt
c+8RTKftzF2P62SU31SLHlRHYt3qQgLcd3zCXZcpCEAxYmcHP8a3TvsdqYaV6z1xrtmflMgkA6Oq
/IaycAwu8BcOgiwEMyDFVJlS7iZMcGHGqbzMJCcqJysDkFFxZ3YH53wFPKD8n1cBLWPI6Gu/6fTT
UKUVmFfeGzZBpwc1n9icQJVlDaH8qq3y9p4GttCgJ3MzOkoAd5pR0dOaqaZ4jOz7sX9xB0DwYcYU
T1lrSI7adkOieebeOWE6Y5XEfGA3NWmJIygKwET6R8u6vkxzXIHZga8fHouXoTNexZnwKwaTeznd
sWzUdZZ954XKx74cf+FgU9d3pnlYCVtuAmahMbKKcJSsXLsN1z05xQjrNMRDb/kqHC/uE8ssZInX
TBdva0L+Jesz1jN0R0OzauS1j2PxM3/wSqrA83lE4Mlzwieg3gSz5/lcSbmPIQU+XJLjUD7HhQO3
ZP9Pnu/GM3wUdDnB6zH3wMnAZ/wDoE71NENIVa8M5TL2TLNQF+RPhIK62MYw1sAS0L5Nn+XNc55d
DfrPoQne9irYDMsEPF06DgZYTJE66ywOTi78Paaq7nh4vGqm4W/p/V6hGJutvGmDugjeHI+a8C2p
3C57Ti21DZXAflwRKHzaGJ2gtNkziAvn2PB/7DdRCLUslsO2PYrcU/QYt1WOKlKp3jExCtiTKecq
qfRXUtV2BB4MKq/ev2leCd8OLGeqoGtu5JkW/3nqhZfCuLFGrd1XkBf16Vkrzfw721mlVUeWVBdL
y30hig+uC+1dETyLyakbHbXheVB1ZOLmkHibuZUcUY8QWN3D7pkJtLtPWaX5C31vyMNekwXug8Wa
Zd6wjOWDPlbXgLesVLl1FDMvSpebdOvpDucO9AdIOHe7C2OstAkZAHzTtIva8SREA+WGcKf4WKrL
FTG0Hop+jmuSX8bYT8Ptz77F+xqbRwN5w0gFnMezqpwjLDg24VZgrhEJbG8tBqpklFowzIKlGaw+
SIYvopORNkCRJWnpP6LM5j8u0e22kzLirLuVvuUCavNC3mv69nMz31IRmwXzTa26KWOzdDyXKoLd
a9mL5hUPGQKKB3GwNio8Hn3g9X7m/860ie4Ki1g4EyXp8m0JEkuNPkUsdlzEwQCzsLyxx0YHwzvk
cyuPjaMq4KE/UKEhsoHNdrMRdW7r/I2TM1AjnfhdjvGR1WMkGG94grhBnGEr83GFN06pAQJfoosy
Jh3Kx77JxQ1Zw8piSjJB3ygi6abpKcJ430CTsZjOwrKPZpO76E6hSuzJfssUuPZvkecK1ly+nD2k
MG7Y8POn1aLGrcWImrCKjqcH3OneQb38IfhTnfg+1++k6JOxKukWBJjYJPI7+qtIszxrrilf+a0a
0iXV8Dsv5+acPjSH8pHJjcm5Xgd1sgy/YWPLMmYo8q0Yh+IkuWkPGlsxzKQ0k87tQlrdmuWdYgkg
MuPb19Gh5hWoYt5Nzirc9QFzho/S0jWIONPc5fTOiAoooc6ZkD28liucwzX0BNxMqddFz90oRI49
D537MzFOEPpbqCV8yVeSkNcutRaCaWIZ+41CKfDKms8hagwqpV+qG+KzBnZz7WQxYQMTjLTr+MOF
B9/8rsOLQCWnDjxAiEgJp/nZ7xCb2AWwVJaiWU70d3sSuRdp7WBiTxh6AzpmcEC2TjODldjdFv1O
NjXqOGJ/1Ox5LfHnpnKYf72f3Josa2Dt4YIr1jEhjk/fvZ7uWTTC+HEdeTzfUBoflNRcNRQ5zZIF
IVnNPk28+6WmGFX/BE4/1q6aGd+gXzTGFcC0nJIp7e65I6+ETjOq+YHwezxyIlNT58YySBYnIYkY
2CcHtqR7KC6jgbjf7Qflwg0+KWobC+2RJyYIffRMQcBo8aEvBLvilEsAzzddnBK9wVzUwLGfGDw5
DZRZCokYktuhzVorWklrIQpRizfNt38etWtPuezKI9dFXe42mq6834V0DWfzYUocOANZoSclNQi5
JMPSiqDTHSJ76MaIhYeTM9X0JiVXJzzPQS+qhZMrYoJlxPmU30tdXNC6u0l9zUioNCsZ0IiEJi4u
97tEcsQRy8wfQ6afkZqgMcEQDrdk5VyUFu34oS8n7+To3buF8BCvbSe9IlELcI1I/d4uoJDgVI17
wJJe1s/u5ob/DCjFYMqHksWn+Py4gZhgFPF2HH9XniiuOFfWZw7ekOQv7z81v/eGv0vtxfSIfaM3
k3RgFiK4MuQbeFbqWrCBJmYx38b13B14a+Y0gAZTxi6iJEUBiqmo4WvxekgrPrXykPxpVUv3ObWr
TCe09Rvtm1Mzsz4QH3933ES82+ZlsEJ3fAGW+DtheQFtSkxfXZAbynb3reci9uMz8Uowb/EdBxjU
QZw4sZk0lovl91jVLmPcbylxKce+m7xAJGD5Sr80PSJ4v1paVVGR41jUmkC4sA4JJlNZ3QSI/v4L
RM4V3lQJoH0Ltvra0OlicJGXZ9a/e1GpL8vQsrpa3a9ZaE09KRirRTlvv70qqXLlUjLVi/s4Cnsh
ogg496qfn/aAkelNr8l/gSIRh55xORuoDf6Xy0lqGKDOuHrI0YAKoRMNRqiX8cFrAfklcl1dBSfW
lZNsS4GS45/RFxrLca2Kqot2Vu45CJmJwohjcYGst2RievxFvSDtU54F6gfFjpIvQKzXPCT91HO2
+x0EpMT0j80W+hqWCiRkL2ARo50msNgaNDK+mnGx1ok6tcGpdin1otpnZIiSjMRK5A0ciIt5z2A7
92aDks5PfpzB7+HnvAwq55Zn3iuA7mH8sPsvC4Vnn8dCbpsof0T/IiRJLQENkC/rOKt7jq1KMxQy
EP+KR/QcHEoS3FZpa13jcO1/1gRzPEn9Jv6b+/AH/OrCzJgZ9qFTmrfvT9ULce7VJ1cPKik42gex
/2r/bXJQzIwepUiJ0DXSZw8APPJgCqxNgHtiPRd+1d4o2MRFAUIv1HPPYHmqlGbiHZXuCaGk4mM4
nGS5C+ZtC/vzbObvd57mQ84Hq4I8h8sSxQ0DknBiUUC04nFfNHTS8D6vPQvl9eWBD2hgDwuQVg+y
ZvV6BYk9mVdQEFW+Tad0zWNAybn/QY9ZcMyvpOjXggnqW4+GTPORSuu//5HsqzVvL4zBNADmlL7Y
yuwKNXVRYSj5rHeQIzArroYp6IP6prMVhO7vEa0qv2ZIfiDWIgv3UdPGGSQ6ccsuLuodt299c9gD
fLybLWFQOCLYkuNN7bOFQDX4jYAM7fF8O7wsNxkPabc4fYJBswzZr/xNTJZX99DwyMP5pbE7msdP
Lg4jIpeJwFVNLHvODOykIKRi1hskeMaz6yKElm10Z7m6lG4VRkmgsCXoR5uhDT4BgJJbyLB0SYH9
xtzQBmp2X8hF+PUrEH0C0HxTOq0LBkpxx5CXNPeBBD6aEb3sdRSMhKLLGKaETo47skQN2fAQqMhT
TdkXMolLqqKhp7Pc0aqEPv3rW+CxGdebIHzVhuH/J9BAZLUBfx63lqgt86G5MsCsBtTPmYHN27nl
k8xnXLX0OOGMtv4P0P1XKlFuV4YBDyIYgVdDrQe37hskdAeOtKWJ/vxvalkLBWCc7/LYOpiyJJ1g
KCLQNgw45bBMV3pyROXJfLoS63j9baemAPW5Gu0q12aojVEKugwA7LnQBDvTRkn3imdHrhefg0Nl
F7QlUGy/DKyVMJEFAa2zUp1xH2RT3WQysQPCqp4n8/5BkyYfifwWbCoW+v5EGv6K6c+W6lHpTOxJ
3fU0K/SifKERxSVkNO9Q72A/N2UXU1409SbbfKSwYvpNN8UDKwv5uO4KhaFQIrTGiwpHtlwRj24j
YJpFi0QcVe3JfDNkP0Yu38BcznFO3zP9Fol65gy4Q+51mOd9bIxW7nQzHrR2JwxM2C34G35sw/dL
p1DYdDFa6fhD4/IHrExZ/YvND2V3Pbvmbqy/aPdDCsaePi33/b+BhKBDUOqfMRLkLvoFq3fMdAlC
0qkmdSNsIG/HH9KUcJqIr5hwh473NRAah7K1IoaPbRmxdW/E1UaMT7RTyQOWl7aTc0rohTZ6jU72
4rM0otrkIFlc8E6e8QaBqJwo11RPrHWjc0eWubtrFoFwVq6n3PlBUBUO0qaHZTsXy9lwUIRK2W8T
7DqT/4qAgC48YFPyKpmRBkyP3K2YZ25cBZJA2TRTQGYWeaAOW3LyfsHR1S5r8nJQO/zD2fDvez4y
V5NZp/yC1KORXHBv1iE8EWLpLzTuaHEbGqpmlpbtElrXiys5bLuI2KGgUek3kRaj6fF6TfLi3WA/
BllM7PUXTsN6ECPnfrLzsMT4GKJMYE+ifbZT+AJ6jrgjMB4ICDx4iVdJt4kn4Sy2XFB0F9dC1/Vg
5QupB/iIxfzMWxC6bljUUS617ljO1dVaAv/4loijCKMMcm5juhKlm/S7Ab0nkvFbu8yxUgQXQ370
kamIgCMXhfljXI+ah9gOrSy2HbrmShh31KnEIlNg2iTq3vdIcV/obQ+Uta7PJnoZ2vk+lVIMiVyR
prc4/iu5GbxDr3U8Tx4S29XhXE/OAJ7kefAB90sAYPmoOXmVLJR5s3nY/o7FgOA0pP6KZ5KuZdZq
yD989i9LHlYI3YdAhTKURy55GAZ1WMpCO/6yFpB1VUM9+s6WSsTZ/YT7twNJVnHgcV5xhSS8PzfW
iglehzNcL0wku7t4lJlPJadm5hpzZzCAfU+NNhSW/CAPxya8pjYplSu/TPHxFdop2apjdtZxwwJ6
5W0A1ncwYiVl65bTO+DU8aG3rmLglwIxiqdWb838C16HkGHKjY3QcBu6/8bvOSMJqM4TcTm1so71
SH2PKwA4CM3ijh1/DJVHUOQMEGOikx0vemq/0aoGY87jfxgzBpvJ4u/9y1Lxp7ZvYLKcBD/J1l/m
iDWnc7wkeRDVVZpVDqtNTeevE86r9/DPOILpt6fVIJroFJ7JWOO5b1pwbwUBWop0YHnBgH8J/xz2
8YnWxSUMc6+8TktDeKiVXEaCkdrbcyKSGN4PRe9M2nKIeu3B42EUX9ft0EicR1IXDHMX27KFhBxv
Xgbu+ek8tmE/MApYDBFjmJ3RWTuIIcMRTEa/+ch2ZkEYB+C/lM3TsuSEk63B4ExlyxcSXj2CPH2U
mQqD4O+744/mmKVO4enq+ZsDy4OsTlnXa+PMIKLTRl4DS+g4E/YNb37ZYeHIomxOLDzywhTxc4N0
e2XX472iBQmkAszXnWnZVSUpG4JwYH17ctt4EyDMk+JFVHodHxpdLp2E81PhXNm2DvFuxRtRGxQY
SIOFtliFJuPsI5csFz18kxUYkC20+VsiXuHRZqspt64o4q+wIes+vBX+0cNBVqPeoai8qdusdeTE
V6yFKS9JLkcxJnQAhU6FOsTKmy7c1RT4n6Yf8iItMzrqS377TNclgyMFS3+Be3OsBaBtRYDDI5kJ
jFPxPxIEND+Qdt4LwwA9E6PCRX/2I0jeLOW4/sI89dCqh9DXouYbpMcHy5eu/htW3UhFDtz0IXzq
6iLPpbrFZL7m+UX2ECQjoi34WofCgjnq8mZo+TYrlOwCbUqxbGax/QVUzim12BKNUhJ7z/53RPaF
P74nI4r9Cf6npTlLvxFhEPe/HAqO57qluGMUwKksc3suMhh7A3YDr7Py5tWJGiJA7PfWYjxkFlTm
EPech3I0dFurv5kb1jdHugP2dp1ozjx1WgDbwnTth8u38ZV4Pz9iWLpj8mIBA9Gz/PYCWBiqpsLR
s7G54TrJjFMVOi3o60MuQuGx9KtIr+5aoNwkB6vv+CiWgqXkovGi0y/Ua+iJudyLMZ4RoX9d60T0
KXIRYcCXuQRxvA/p+bH6bs1ziAz0UR3mAV3Y66+DKqhVb9VT4nwstbNsLmEjF/aG6kuRjPx82qio
5GQO5zq76ln57wBFJoHvfjOGnQobbqB5AgZ1GI8Voh2JAuSQOr+szrhpJgYZJFg2VGDboWezDEOo
bAl/tnLlb2dm9xZT1xu4gAZGv4L/wuSKi0nOg+dvngmy8+AaYqacGICVsLjiyNftI/mDiC/A/Cls
+8foZEEgIQ30+bKSdPijHJe8tcdGk0d1AtHcGwyja/QxHoZ31FjTk8YAmoMRiTcOGl72meSNjoIk
HjCcRLCx/4QmCR+M+CBo9xvhfRJqM51HYEp2nMh1pRYmcUQ+SEfVOzpTUP3Mgnso7x4bC7r03YeO
QqxQpYc5YuFQSiqybq4NeP9XfSQlyUyP5bsmOl9l4kLrZAf1JSOFCC7VoNtz54pHHcc+O57pl7Lh
dRJ4xhmYLJCKNAJuUCYP+TdW5l+BFqbOL/oYmt58bb/NIe3yybcxq57Cg4+azvzHDlM17yErt6g5
EtRqHkvwCUO50Q5WigB0VHpDgvl+lZCNovn8hz2lhIk5GJsoHY0hyQsn2/1vnIjyajtTooocA2qw
ksY4vUkciWzLqSM6Caoizb/wTjt0i6YNRg3HgqQHIRqJGt7T7KD7/7puSwuoQvsae/KkHHs2iyVK
BHqy7m3/J2OABOfC1Hsxy1BJR3Cp5vb44G4fVKPQ+sSjmPCHZb7jzEirl/qqlUbMf08brbn0Jh4A
foTYX/6c26bJvXWGDjD+x+qS8FHbcmUZnm7gnV/2kBF3D9ZZOgsuqs7qIkL0Sn5Mq9nLpESSwVSh
NjuR9xbGrqhMa6b4s5WGJiHetLfFQng+BqvSb1+kF0YSHV6pYV8ZiDPGsUeOqu01gD5R5kxPFiy5
X16HlQijcFomAr8uJh4dbi6ELfpucyBxXf3qV++EiKKm8zXePSdOvcS4nWHH/NlnTwM8Jw3/faOV
F7eLHFgnCubSNtMOL9Fasg3le+QgxToPGPThEuZ9sdgzh4bhN6c4H6E4TXcbEo1hx0n/RAWHfQUm
Tfs6ghgMWT0wBQRIFTNzWTjhpWRawUID5Rssef/HKGLBlxcIMDk89XUzQRFC5ZTxdmn9TlwKfOho
Q2BE62ah4UaQ1n39mAA4CKE2M+dRBUxix7/+RmHbo8dK6B8L33SaMrzsC8ixQjs8xBslwh7fuchI
Sl5/q4zder2dYTsdeDhelh4wCC3pvSX1gq03NZfFkBlZIHLs5zFuxK0zrpBw8WYitDtk+dqLWLtS
DBGqlPxtWG4A5eWGm0XH8aOdsnENELT1wMiTpfFaXjVuizAlAVcvr4L16cfVRxnLDGgwnhVcTWZ4
QDLWt3C/DRQCuVN20Z1Km++tsNkInuBZT5Qsfi43Mx2K/qQ+dUulHMs6u0/0m/yaSJ5teeKpqNlV
GemZUVk3awp60sHKYsPXkGErFmeaeRb1bvftU4qzmXY4diWsGZt8cxJwuUTJOZisMx0WGfTFBtAw
58Ln/0OlsHvtfrddjxRQJv/bYR9pPNXeduNzM6fc/OJ4RAB1rSlmssgV+Wo98BCBR7Q/JK459fzD
XPqY/pcf/EwN1m644ElPbvyD9MAwilzKFwQGvu8lOKTFX61CDf/QxDrVF4TnN74ineTiPyo7jlh6
f2AOTRkWdu/uIQcO5ECxXB7JJZC0ge3KZfnRxkb4aOxqNVuBu8n/PE1gq4uS0RAsRYCmQSCdupot
9lEqrPD8piqtuf1iSLBrzuz785/CuCsq1M4YXUMH9WvpnCclSWVTJLvgsMjigGgtPy5SBCsxfUZw
WRlfhU0fBOu2r0gDwIw6no5w0PziLnSbsXYCFF1MuXAByhJRrTm8XtitjrOoyK+cfNN9WS9VC/KJ
uwOakBEGmT31/FFjCTw0oP2VOsi0GiISHWnOcvopDTYHKXne5egdLP8ZrdeYBeEyFyOCrmz5aOiK
ICNp2/83PE6SIGLdkfPr3v+eMRJZAqFw1MRQe2zi9SXtOM3KREJVCwOMz3PrmC4NTThcHoDlOUSY
9oIrVuSuE9KnHM6IB9sX4Wojv45n6NXD6JKozjkyOBI46bGml3mPVlwtybVhTkmJ2OGI/VhMJ6LW
gdQymqaRbWJbUyP2PuxCCRwfB81YChmqzMA4SWuxhq8XQE8HuxtPjqRwGuD8xaNtPhGM1PMvn2BQ
UhEEQyBpGtcxXIH52q3ZDI0UF/ZICwhYeq/3tDgNwNg2SRBEmCBxyQEyQecxOvwAYfMKsCSpJiFR
IpvRHzExB5cK9dpSnCzmp4w2Q1jN0bmvS1hfHteZEHeJwuQUObcCG/js0Hk+jp4+Ut/p+Auen3RH
wA3+NUG3K8BqmT036f/AIyYNR8P9hK837GIdin2Ll5JqSF1wLt9694ydQH2eDW5ZSt/1zNxfYSL4
ERiW+wTT0NmpkczmbrlNC11xpRWtup8+CmExPWgVW31Co16Pgp+5ETYG5jkfbhzBcG2VCFRFGqPQ
dzeF8vu+EzxxRQBAi95OOo8zxxBeC6aCpXkGkC6y4C3LlJB5cdtvJuWknOb8E3/c4FEGidJH/9RF
9co40y3AjsMRqKAuOm1lSQ5UtnRyf18OTcrbcI2n0kd1NBj3BuZiGl7Y6qpKvwfRq0X7isWzl1hs
WKaKG50obOiSoDdfvpmDRc7FyTa/fgRctjszu1OKllHSwXiw3SH7UxMSaZ3aoezg9bkZiLdiX2mZ
6pavA/RXUCILWB7Gw5rRh8TQAMPknNGOA8zoT4y2aNdN4zNHUE23S0FBuHDCOa+E6ZQHLwl1uT1M
Jm8hI5/EXzFVVF29rQ/UhpuENcUpPj3eHKDDm5mX+I01nINiMjOmR1Lq6aYnt3B54EUNH7EcFRNV
3WrpygHYUUbJeTqgnjGVvrG0g0fJMM0CzYGO1rnt
`protect end_protected
