`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eKWOI6UNAzTyoMOd5jT5prexud1j7tO7RWxjl7uw+BChyG5RovhckwXUF3eTW2W+sbM+Lmu6noKZ
7lYZaVSi3Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GYc8oMs4Jyqcf37EkXIDqE/YS/dsXOir1P+2yuTZVP0f7++IsAgNMhE4jQ02ziHHLy5cjMEVQOcp
ubTjGNvG5opiW9eb4EaToiN8x85O5GJKlCRIXeBXKVyvcT/tF9lTLdlm5mn+JllnnGaflG59MMg7
UVoisyk/bMQf43rV61g=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ncj494a6N9Fuj1Fd0e3HapquRQnqubEzA+P5GnfVo3gXJ9FYUGijv2c11cIhchrXLwvntGQRNcx5
XEtYoVEJYnUewEPK3tuqb5KoVQH0PUMMjlPkZypnqtEyjv4ArwLaYb9HlWtqz/rKLBpbdgMV06rH
inDfqds5zfaKY73NjX2uNP32fb3DqMxYTL50uPWZk36fdJWRNfTdK/wIt8PKdzt7SfxrA6gPgZAM
nZW7qKZEGVDBST1SsBDHq3/VpjdYapXGkLm5Pevg2UjRmEAIeJc1Uf9d0iPFaXLcqzmkCzhLT0Ju
bSgRp8SVAJX3f4hyHQRI4L8RkAIUGrVs+5fiSw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
OcHqOzyrH4rO/VGvg+DXlvViOxYOO1yKdYOXzVjprFaTWJ+kU2JYKYRijKDcOakcRkzxZNbpAifN
J7a8H56ExXBG/6K1yuBScwln4vsFqf8NZIBLU8vzqujDTXpTxuekD5cUi+bXLRdbXoPulckp+45q
/z0O/cJWNYAR87sGJ1c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pGak0Ax4Irit9h2RpEorUU8qF4PYohRLpwH0ewoWu77u9RttYNa9Klc5zuseyqzXzboB/iHWtvE1
Raqgh9Yhr8csgoZ1h/GoyWnvJgjA20e5Bmb99kmaE1MdjFXLv/nYMbU+Xt87Z9uA/1vPwZVGeags
TZh0gSeuyJ6Oj9DWiYY74F2dbek6SfNHzrJVxnWkJPWbW5CClSxBcZYxFBiWW8xqHU9h7rkKNtuh
LdJCfePtrPS9E6WKn/zvTJplKegnsaytZO2Oo3T4uGzjxquTOix2ZVmY3XVPfO2Phi4Rk0xZwuEN
j9lKHsyO5/2LqPTRL1PmdEjEbYAtxz/tNd0e/w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6848)
`protect data_block
F+p/csokcgE5WVJMEIYPOL4kwg5JYr40jvtv/lsl4GqtfujbgO7vZcTpI3OCagPNC0Lr1jigmSsf
cP2mDbhXpOHo8JdU/wSQsMeJG24C8xoPSKaYXHwyOalpbGLB50p2g+0aHqK3qcIcwLa8wMxyWs3s
E7Alx0t5qY0nSsIt/eRZMLk0W16bb+mlnELtcMVXiADLua1ZtTjNoAzDYl+xOdvzyPoZlz+732da
JAOfvF4svtKExKjB4BzJR/m6ok//wzeAlCW5xitk/2NhEe975K9Az7J+MnTJR0zE3dgRClmGEHQn
fFL7JTpOx2Nt1NI08OMUgH9bqj3DWxntcNY7FchtjrT3b3Ku8MOtE6wkxRyvbPhOxcic9L6PCnQI
FJR8hd3PsDXrruiV19QrLEYYntI3XO4KRF7hH19/awHHkdtru6gTY22oHlyv1Y7mRmWWwVD3njZ+
FaxsAfSR1gqMXEG7HRHYLFhUdn5qHVouSQ83UDh8gg5Pk0mgu90ttDYkCQHPwb3HPNUz6JpFHfTQ
Gc7kZbKzLNFgukhnvp8fyX9AfRRyhIhEcNQMDjVCsRCKmFBTozvXavsX3/cBDShUPOTYfve3k8Xf
URr1yeNQEnZwsmS+7wR7Ix/sAllU2eieFnN6S0edwF2x1seUZ4FvnSPaNPyVPpd1h+XPJjADDcd2
tTPrRT8M4Jlrn3Y/pRAknAtmFLytqwU4ij2BYGhfCc81XIYKoa3r9GUjHNqNyt3ZZC61rJnbKC/R
zt4HmL3EUCb2Jsh0ydvwJL+4he0dqs40NAP88KJiGy6dVP66YYt0Z15HQg8mL1ZUwSg1BrpNL74+
7c3kNulKy0bDLCc9bZNF5zVWlZJAXN4AdgQ4uYHq2ubgXMrH5a7FIS+95FFqgPL41pjPxn/fBx2h
YRosU57UISgeXlDLDwbCz7pia/gWvx4TQ7aFiiXI87vBh5T4ZWZGa6Lbdhxe96OUXjwEmtqj2tfG
I3P6p7KgXFTVQcNx5TEceUJuZDXzVrbHJJflNGN7SaNgMJLOi9JnWCjyc/egm0m2jsOuiXgtHfmJ
9h0Lh+I3mhayLEQ42jtSZwNpICak+oFrYHutvqgNRFVBBT+tO7J9vesBVfbScmHj7WqVgT8gGHlc
Th7LtYNPljYp2UIDXHoKZBpZy8lv4qpvbGKiJG+NWmi2LAvZGPKCZtgiOmpgrRmzZvzYXlRl0N8n
SW3Zm4fqp9xp9jkXYbaqCVOwltX3y4wpj4PNI/XldgwLlHxsgDUTdXZWjfkeUHEBsxQV/GHk1a5z
5AoO7GDIxQPu4fGSLT5YuqT00Y7Zbcz6dsYzkllW1Ln7PBs13XMRUdV/sbWRvEDayCljDyT5bhfO
cY481L1kfrWOxbDW63ZGeoDMdQczYlowBQrb6lH9C9WgrfN1iF27kU8Xg6N+0MTlb/n3WdBIz1Af
iTfrHUpot/eF3gnXeP2Iyn8+OypL8Oqd+VhKJeCd5vCJUykdgm147rOpf/lHaP/Dvo5mBpLgZQpc
1Zbm+7YCRRzx/CILkjVACCS+DaZvXt51CJsR+M0OYPduCHFyinwP1dDk3y/URBVFuSGLDsrIDr2t
zcsVSK7zZJxORb6zHoehpkXolYs5/B1hhAzsMxWaSmc31UZsu12T5874/Lm+GjC+khYSjTGrX1iA
bVV2NkREP8kd6r4pgfNavTcFd/95lgy0Ca5OpkA0yGA/F4yq9XOhIKf6xKsc/YKFO3on+MHxVBVZ
GBS/3ysqWO8jdu7y45/7TIaEg5ueV4k0VrBwPEA0Cvq5fTnWxUiobpDFE2T9nK6XFYE2FlLgjzS9
zIWSc3lzM12T9YhJ/Ywpi8l8OCU/YOX4qKtZUMv+CQTmuKhegmSfnSv93G6O8TjDi+GA38XAaYdF
tcC5JJ0XqHaSdaAmxAPUwnLDNlqrlb7O6j2vfmcr0yMWYMZCaIFXDRIaWMS/YJhgJqEQry8LgW39
nSmsG9R621IVTXoWuHoL/G4cI27spazOvN2TVCD7FCd4sxtujfWcDdThzCPOtrWo+EHolQlLTXuH
z+eJz4Vz8c7kuBccuiSB21DyOhnwv7LJTdAuYNqY1HPIYeOpQLHytqh1zdY8Brxh7n3pg5VKxfQs
oiqKNTZ/9nSp7iwKgKFDLXVcDLheAbtRjWWG49X44ovGUpPlVt6xEDxpZTEhtQ2Qs9q6rMs/jj9e
zCl8Ucewu2iYna0ujmsa8Bucglx1T5ftgYEKpEpeMh+5T9t0U+RLXc4bHcf6gkmkOkZ9BFtLWudZ
wkv3ocPHMXpjovdOatOanNcraekmiO/dIovCC2/O2k4gJ43Ca5YjfcffNv05+FMzzeO2L61tKV/4
rHMbhNAcO1yA538qznS8Qar8ijJbtsGGjeuNmqJ5k5P+fw+1EMljdFYCLFnLMe0+ftFvHXo2SUUn
AOjxSVz+KtG7SN0taQYfvDDrjzgP5tva3/JjlH6WCx3lOhrTf07bNYHkeU7YbPtyCxMoSubka9p7
ceuuDNGPvuQXLD5mfPUY5M4Pr1KYwrma/dhv2sQVGzYLJNbhRVqTUeXG2Duq8JwNKT7WMPfxQ0RW
DCgYwzVapfLU8oNSVAV2nv6X16CjiJ0QB+XnNsoquzulJ5EdJevawA4UJ+meyPplOYQWEb11SZ0P
PUjJPcWMpFk2jp3ekryUQawnHSWBt/Jolt6CeYlJ/sZjZxKo8A2eiJSqibFN7HBU9yUXDbH+MBYi
pQ6LtLQFYAqER6HgjKFoAEiNj5wSGw/xpqn9ZzwDKdg9hXlgHqfIivIxSts4aRalzDhR8Ii1Ljsj
wkFjnfNCD/uV416FsmLNJ5ND5GfZvGHgHqFU7YPrTRvDsfGyg9EkDKygv2zIbv4XL6UNyITuA9IL
E9c5WZtls9WoIF3xWswQf5bj/TlgqPVN6dlzevrFV51dpKt9elfebSNCriEQH/btZoexlQKzwxwM
seKJ3vX8sVOpaUY2YS0bP6vk6zK98iWve7z8g/JKJS3dxfMsj0eYtbttKdwptfy5MbRuBmunQqhu
NgQSCbC4drGMof4d9msxzSOPO7Dd31iqWjoHIUzgva64LJDk1VIxth0g10/RrJyzrxu31Pzm7h8X
Sxm/lpEp9RQOrG7yXL8ATHVZ0NvxgC3gZghZfc/PvCm+UxgjSZgz+/l0fFWEqz73si+Lr+Ht9+ie
87NPfCUVf0jrKEiuHbeQ+nRXMm6xCCzeSc9aI9L6HdKacMgy09nvbP1sr1qpMGb8+qKsyKpu4aRK
i4WlymjiSKt+Kwm3D+IpI4CLUU2Ykoe8hknjkHvbVoftL7eEJj+HFe02KYXBxVGlje8aAEAVAaj9
BrA1J4F2cH4h3RnafvpLpLyOM1CHL+37vs2G7kWTC+sQyso1SVAPtw63ccUzvbhHnnRSozAGZSs7
FTLW1phm87HoRF4MaUCYojyLhyJj/6cujw+TeqrCSfl8zfZa2l76bGkEPB9vUADo5WghPqud7sBX
C8cWbQ9MIznZPZmTJ9Q8TUpIOiKuSPFjN9infJi/W3GNyoMXfFVHvlLwVhTdKRVB+hSFhmp91Kn1
M70Idl2j5dlKSRJS/Nd/0PrEe3nc2USY71bQvBHbU39yd2oi16NsI2x2WGzuoVEza9pUpHHkeXSG
kV47bk+U9q7PZlFraIZ/gR9dw47XEvEPaN/xnFIzR0LN0/vnlmhG+HG8qmKpUrm4kjHxmYk0wU0b
eXj/Uuf4b4d4WjrCYjBGag1/s01Fyu1Cy6EWjWHKaOS+GFwPm7JHk+HuCHXKWdqyQ7N9hWZfIbwh
PIVutq/d25zUIPi+jRFKsLjQIQsUceZ7SUakzjb8OxGOFKELxC1P7un4/e8TTA53J0ls+0PFZqIC
q7UPIJkdbEJA3uBrV/TZOTYDnYYGs6scn7QvetcPkQhLjThDEDm+CaGsQpIEvtIrRNxenxz05kkZ
aBAf4m/cEwHM1CYRHkJUTpQ+cPC1WkA6+yMLw1LoD8zdygcynguibb1soOTJLvKURqFS1Fucx/bJ
dKtfZv/SWGY7xvSXqEfUNUUJRqOmIF1PSuYXiqM1C1wufv+3h2Zv4/Vl7AJgWFTYvjiG+rOk0V3c
iRKql1GCoA778c5HaoR/rLw8Q7pJ6mRDwChXR4iyYLCPugBxO0ZXYwCKLWlx5m8RUPG966ICbFVT
Uu/VFJcA/6UdCbAYvcCpjr/HIKPfD7y26j2x1nOkFbGkfuSa14Dn/wb6moaOgsnp1/tQCA6aizOV
qrGitSaFvEE24g4ETp57FaWZra5RfKpIL9Ah0SG4ZoC6mEGesjsO1fSf+TyCAFY30y/+RVHiaUF4
v6U0UTnTq62nZGa8cPqhgOyYbqzw1yT48GlN0zUOmpeV90DCqzO4zgM387KY32opNTSpHCEKMR7S
hjjl8WTzxbIP/glvp5z9YtFVgt5ONChgA3R+AjX/0mZ0CDLoFhfkpKKDhhG5Hcma9MMrfltixDm3
6z3rd8QDYPxRJ1RgzZofHidtFz7H+DyiAhdOpUyKz6QXAQGlvmiRa7598iyDnJu2ym8mzTgQdMTk
I2pFlxR72Jy9U/9pWE4BYMUmK5g2riGzz4ZJMqj10N5HVTxDKbC7EJ2HLjw+gePXHwvxoxKC1qgB
zUFylXS+Cv8wiKv1swQvyDNKAvcMjxnVEahxjtcxvnExbOKS4LEZn/o0fcSZvSquzTLVeMQpA631
1spYajWzk6pmrZc6wDC8rFaCM/6TOG2ikbPkCLReWxPImJEwK/c/sTMGwbb4f+k3x3Es9G5oswhf
GZKA09ktIAgnweKC4tk1RTjhkVf9piC2c0FfbgFY6AiRl1ZzMAuf6oPWme8xa7uVtyOkgx9Wt521
BQgaehRh1hdygOtMMQiVmLk3OJiNZFrF2K/dl8JR3e9sUaSJiMSDyxKQ/wiIlwm7zNnliBN7pTAS
cUoW+W3dXriNy8HgDVQMqE9/PFB2fxGNBRVkLnJlDpf9HTq2CwGi4XwowmrGjx3SzzeKeU+q+gfG
ypuRZHeI10bIVpIcJ3wORAWZRBt0a2MwzkM4qcj7cMo0MK+2E/pXSvo68rlMno2wVIr4LmfYrtb8
/IppzIp4bGsAyYAdW3zNzS6pDAFadtoY0E33bJWDH6GsL9jSEdV+4Tx5PMdU4MjalgiJdVgNxXtM
y5UPD5y/0Cpmgs0zNYgaVA3isjTHmekjYW3Dtw0Dyyr5p2x1160gtwDtW+ao6ONNsqJp9a7AbwxV
Wy81G+CtApcqa0pKDV0G1tvdWOERoMGQI9/+fOs9f/5IL5y8Tgp7175cDhEwps4UZJFAR8Pf67VA
yoHFKzeGqiRhDslGCPaCKwgkprNz96+AnCUSiTwZFrM3020jENO2O+4M+H9nKaDKgUPYxcsu6Xxm
cbLtnI6X0k8ymN/epJdkFmYlsqyOuOIvqN6/e/oon7dKr+H7XNjfb1xnmtJr7Pwuxemt969CgllJ
4trLXIJGoagX7Ss+jh7XxaKkcOdf+xaoFQn3F1C/IUD1hnkg5swzdPKkYFyXX5naoEmSDN3MQ9VY
eMEyWe4NemjnPsZnL5yztq1r8rzYhgMKiHyFEb5JhXWmekGpY0Aaoklu7KkWrgUecvajoiBtXwU5
qgFetpYQ7zxlq46nDxSvQJC5Yk+4b8Cg5O/FUfvtQ8l8eo3iSAJtHws6AXukYjICp8gxsxcYeQgM
b62EebqRm3/dB3grZUW7SdVdEbrXSVOSP9EC1Qdj0wpQlFcYUHBs6ufKLiHJqkTj9QxFWMA33WgU
IHd8MT/UukP7YyT9Cc6/BhXkJGssx4wWJg9PzV4pNXVsJb5XM9JSb4KXGo9kwsRzEv0wisbKFn9d
CONAuRKy6j8eX6I0UufSyFHbZuZWbNMYh3+C4X4W+1U4UkfwLFTslD3QS19WsSLqPB8mgE9729nH
zAv52pzV2GXyElJm3mrWLfN48rWrL7fLBe7v35RIckTQIhf4kFrpqeRdhcG+sJ4sbSsFksFfb5ng
PFeHwKNLwkxAisY58QVDx6Yj+QDVdI88zcjiyDKd+MjF27OPsHuKTNWtoTefZ+x16+R7M+WpVOKS
KL9pYqLO/PCnICnOfd1Ofcl9D2xbQkas4zbvPMV/ksSgPTM5rCxx6M/TbYw4QUjRmCOTXuPNUAVs
N/Rd6lCcFedKeZ/qNjJvHd2mLeX9bOA/UYojtid7s9KiFOWFHTipffD46NIgdQKDZeqqkwHj6QS5
D7yYD5/LgZqMXFwYuSPQOPJJ8HM6QPYD2IWPX16Z/LamXeyLWjfl1KIx4Xe//Nu4fV+nbfSYbyza
l10F3A/crbiQaPZXJGBgTcTJsB0S39x+/aMPEFCsHgXEkYQnlr9pbsXbvcWMwY1YacScSr4ryE26
q8xuFqSvQ0f2kBR2lTaekbNLLVrQ9dVqmDAvVedRCaVG4X4pyyJ2qDNxdq/z208hmbrhSafNCVge
/4sNB1Gp2CzCCddd5W9/WnfTCcPZHdfnHZnpkChAh+oXB9IJDC0cGpPCQroRdC/SDyrNFbZc/oSR
VsAZh46yAUlF9tz2avnMQqopVsJ8FnyJDomnIYJ2T1juUt25cdz/W0LP+nwKBAPUoeb48osB1C2H
RpDeWlr0RuCm4q9K1rRijVrMKJvDceRYp/mVpSWx+vRKyDtthqvIpKjv1CvAs4vJdFJlyPCaVAaS
PWKMIwvf1kF0IzbRNnHo1BxM3on0xQ0jWjJbjYcRBeASd2ToPTrsH9DirRFPZowHgL+JBIJk/yvi
aje4JyeJqOPJYfbnhWv6ff53Cwg+MNLReyjMj+cPfilnY57wnRvo5qGukG43LSt8kLvVgCALvXHL
ggm01tEIPq6PEMkrZ/eW6WJ//16EbsBt6SFGqw7lO7q031h3PPLCt82a4GDAKhxJhC/HV+ZPTuMs
sfb3zLNeqfr+DikVFWcFNGhJ3cYv6V4gJJ+ADlzBdGfth6u9sJ+Cgmv/af1ewYcztZCADEZWznci
k9IFxNm3Iooa2EB6Gn6dQkPV747Zoj91EtxPrD9nbRQK99XI6Y84nR1LkD3osusM87mzigurpZV9
VDFIGane+Be66Jrn3JYjvf3s0FByFlOwZpyQP7Bvp0PSHXP9+6X8+TjFk6/iGhbsN1E8yEy1Unle
ZQWgWTiYndUE494Uw5pMfoN6vnQJ9EtLCXE1aW0LUt4kQm4gLc5SSLAU24Wh/dgWRmMzlJN0jEqD
Zv9HHrfrlZ2bsOMoiUnj+p5xGItS6pEVRXtnhyv1Say6EIsNc4JkuP6C5dbpOElKCvGqpSO+qmwp
FQQdrOahss++lU8yciUx3wnXTmPi7yCZioB3oVy3pDLwSM8WwZ5h1PoGuHfbtknltnTkRgjGpk8y
rxt/o3HWOtkyO6rDPFHZL1328mDbLzPO02kkCq5cj1ZyYbwmlivB3Ofp9FMmwoyEyVONmtRkRcvk
ilSPqWN+WIq1CXdlroBqvL8N4+driAGWkFeKxKgN4CGW6JukzxARen09jHO7SWO+KvpFTwvfIJ/D
45ZLIwt0VchH7xn1jmJL310v8cnL2qI1vMEcHibc2V63gG3sNBDUKLZVLSzEFSvCWgg1wLcAfBLI
PxyTmqE7kDxlKP2WPfJVllGQjhMtyDZ7F5HDKVo19fDQVAwRj+rK2b+pWRLnwXK327TTh1oZmWsh
YyiXQEKrx0DxGJ0Tg0jOmdcpnXnUc8pfCQgHO/F1eGqBLhmuTOc46zv6vle/LXCcPEWxzn0H74q4
FQaTZZCBNxKpKKz+zsBjc9FZov6Tx34tqCrE13nDfRVS7q2D0lU11mt7dfcd5xCZ+zurzCcSzuHk
G+XT6SdVj2VSBt/sRdWrCUlg0NoGH3C+JlfmXsXIgvZpS1Tju8SCdFlXt4C2/H3fy+D2wG8Af5gb
7qDMKK8TVKGOAYtKIG8XN8cXkV+ybj+GngB5ccpguIQ/hZG4D8WM8g3j/qxNvfnsWL7haTUgs3lL
96Py2dzaMdAKhzkzTJ8CWpDYhMSOcSyIYUEqHhowyzUlwXk3SmlKPULhaOXD+7VFlQ1s8K4SvMc8
B+BeJM57fOavXh0UWeGyQirnwW+HxxDfxAQYQWRBH0zJ2m91t/6wmIMRncpWhZGsTsAojamA26w6
9Q0i2iToDy82UN4+flbPIqEYynmS/dC8rfdfvnXF88LOQ8KSlGT6ZatdEoVquAWTRDX/pG2VjP6G
3N+VcR38iuAx82UxElmV3XEeg39UES5UbONd1Fjo7Ei1Hj9a5bMjJGmilalK5f8pkvSXcZ8423jC
oOCni+qSeXvkkzo9ug9rl87F1JHMepnJ2SQbmk8mrlSb/8F2kSy0mMZmPmjfMB5Xh5qEuR8QhcQF
rqTJ38idEYs8CoQC3QAjO+aPACjp8n0+kZnsmpwqisJvQXPK3Vl8hXo5mhp/qhp1WycpuYkhLQft
KTqa9Olmjhz8ME8Rnz/yf+wvd4YkPftwXW1NroOWuh6g/iMs9SB5setU6/FYrzdB80lRdzVmAobU
TYjypugK+tFAo5cPWnHhs/vlBID5sr/VTMDY8+83bGFIPql7Mt1G6HZLigxUz7EKPIbUByY9bPjZ
IrSUMpfUDp5ETIW8YuodohXk52o3dZ+Xf2X9XaemaMz8Eqhnre0+PmS6gVpLzypqyFJdV1YBz1wB
ACmaIzh3UnoCDjMyB5+X07AiGJrrXd+gV6K6p94u57DBjxLmeUhyKkGluSzmR9KsiCfOc7gpKCUM
opKy6lRAxA92eA0tRzHDsQoymZBAfNjCwlw+8LrS/w+V0bqzkM2d/phctf2sNFQhX9odkxezHLkD
Q4fSbJVvNVH6bfe6KtyPknERH0J0mmnBL350ivYt4s2/ZS38u/UiLkBpx1A7xusWhnlzTI7ykkA/
qR/tLVj6YDh07eSob32DzjK6LNKLBO2o5muTGGrMTwwKW4WiqSbIJf4p2z3QgGOPYYqvAX23kOQV
6zc/7JYvaxGbgLXTWxgkvYIJKEY4vZWpZ1AyHhVegWg+xzuwieeTF7BwvX0QPcyCvVRAXaUFsXOD
ObfuzpP5UZU5rp3tL4mO869nwP0XIwkyqKRzQz3/QWrul2lYLth26P9ZV5zlA5WJE2dr7LgXXRmE
ZSyR2de3VIA=
`protect end_protected
