`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fR3mubjMxbTpBXawoQGNg0W6BJxqqNvXErchj2MKo/20shmyfPlKVApRIYIS+n1cekvXMNGRDsVv
fJBrza9Oaw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MUSkvatgybT0vsIGvuarv4pHfjasfOoehAHY11VrE+nBwMH9dUhaNGoNkOYpcA9kWxk8qGxHV0nS
M9q58qDlsNi+pFrWehn+CGwpCT6fw+JhvYks/7pIkhxLkYhWKKr5lmp0YX7knhdhEaW4WFpzz/iW
WY8W2UdskxzhTVe6Grg=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
m1j1yW+q4q6Pdm2biTkP85utoYt9bS6SCniHb7BZtB4MFQaVIlrBEUUap+EF8kUDDOSV1qZ4kVxi
il8uxCI7/qdZRa+0wK1zK2V8MTX5Xobi+JJHCKc4i4+zDVJnU9yI3wNkBjTx4RzRGq/1EgC8uvmI
Bz+GrV3+pKBfy4n9cI5KZ2rHRLM5BKJrN5hWsLWS5T5PoALIVaOh9aA0z+EqWILYDvZIHryks9eG
1iYePZyWv4ZbMFa1FaCIFTnEBNrT0rSfnB2LhFxCC0lDxs9a+3VMxFtbZtLDEj9PznWLtF8P52I+
h83ho3GFtPims61RXiNXZCYL3hWy5lDCvNfVlw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XtlZnIcVmhsDmIcIaLMwluooHhmS01x+64Tn16G2BdFLJLILi3sH0lIt22yrD9jdhEyPw3Wl/g1S
KMFZewBYU3l0WbV9YOhHCDF+3W561JdncMGth8+BrCsLyGiYm69WojC/hZp2dWmhePOYZbSCDaEa
baSBvAWYcCjxU0ekEmk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yo/ZR8z1289CRFS0I5fhYNKb7L4t4sncboYuK5z1p2wK5dcKQVPDberMAAeEht2TNVyE/RoIJyxD
NGJsF14862Ylcoaqi8JgIFjiQup+rhWZsR244dggQdKzFH0JQq9aBOgA5bhz318pDHnhpeiR0inR
VxTWmGXmhNMAZMAx52+Rxi2opn3sFgHcizJXWqJQx4cgPsAR3qLrtAPALLPP2kzmFTzSMiEDI7Q9
6bs4IuVGhG91txI6UYAjCbNkCuD5kVr1GUQ1gXH4eNfe9+CVPC+/kWayifmNIlq+zsF32DkJfDDK
npFw2soGec5Jy7uAvLVLx2zY5+1l+B2vJOx/gA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12224)
`protect data_block
vGpBH/8ieuZ0wkeQWft9zNq0Ikj1XYZoS/iuDc+X+T4LLmqgxZFVl6dn6wiBHWY5AJMhCiXemPxJ
7Ht0Cu+dt8TRHsYuzPCuDZKlsfBQUVkfOQ0TiWq21FLPQA50Q33SeEC9/y4HRELwz0VBvm0D3R4N
O3jBHv5NPY6V/9nGhmMyqH67qGFrmoyZMKrlvY0+xG06oXlHn/4kiUcdWZ9gnQamkm6h75jhztmh
9gG3rytlV2a72VxcfWLz3z8XPZ/qEPAFtU4ZYxeDGhqBFyWtm7SlG+0ArOqQ/RkkytxeofZSRwiy
5HejtVFnzr/orIwLaDqIQIGZoD2gE0iAZZJOfZ2BbEzykqhLwMdGaenCUVX7GsqctLXH3DQeC7N8
yqI4k9mPZzuNh9abxoAHSSbZVH7w7Lq7iV8/M9SsKo8Zsv844HvRfY/1RU5X5FxTVjEmuojLeodS
D4QqU+sIBU8sccpWFBWBZlMAzQMmsrOM9cPcYPVNXVeAw5P2EnjrY5eBouS35peqB9ho1SbPg9zm
532CJyFjF0sS1uSGnXWcUbK2K0PFLCMhwk1shL0RHhxe4hWlQbp2QZ+uOgVvaPfZGqphweB8xsjZ
cY7U1Uqpg6aFUu4FLNrpDvMs+kZEQGnqy1bu4n8yA3q1tPNjKBBeTmqv08EU0CVCK70DM/fvuXvI
TrrJKhZK5QYo4pE2FupQgL+Qq8VsF0AiFhUCOMvvM/1Z2mAzb/WrXqOUgeHF+IO2vEADcW/pCCkO
3O9bMQsYG4YPzMmpWWIoZ+7Zgt8K9kvoCXyCsId6RIvpAZOcVzzP7N25uQuwCc4vJfxjcsjK3ygL
6+5LOTG5Ox7EQr+/6vabVd0tvu8Dp0np4XXHatwB14AFttdMNIiVqoEZ8F/q7bAH7UvaVXlFVWgS
+QAcKN7TqBkf5pUB0LzMb9LdSiNNPQEOfW21t+4UajjTNKOWmV64yHaFszStF28tGgY8sb2aY2Hv
djjIKle+6URt/BMKf4GqUvObwRYfWDN2olub/NnK+RlmPFVyEuwJrmuN201j+NCJdPEPqQiDuOag
ia0mJADOu/kswNvyTHPRErLyPZ+yKWf26o6Bs2EC2FJU9gIK/TWnN2o73F2eN1W94rsXZA//Vn5R
o0gzGlc+3G46S+kB2Bz0XjN7PQ8A+quMP7ban8fZdIJgESo9Uszuw5Jhu6iFKMzUQiNOyAw5/+Z6
fJMVIOHu0RiDuIx3D4Nk/yG1+hWDZuPVQSUargN0J88C+aUismzLjcdBy4eHAXiXITYGBn5XBPZJ
wOEOZIg6kJeHr3GoWn/h0qYNcQVuGJgTq8OTGHww+uL+7z3dgcjwhI4DODGRFvH3VmU65zo5cU/6
WRjJEb3Sprpf6k2c2WXer83uINJyPdDvyFeLrgJfM3BdHWn0Vh4tlZHL7Z+61BdK5mRDdAJ0TXxY
ViqEM7VtuyRREzvFwiajbNW/Xr3h6KjqCtnNzREzTdVUDEk7QqKX1h85eD9Uk6tFHe0tCImPVO70
wqP33dIzYNbovobErNB6Q0ulGAvbG8J0s5dyHb8tKGdjC0glHF98jtjJVWwHad1ualxgRL5p/Kga
f7FdUDPvs7mn70PqJiCzqVHHWynbLTEzxok+Ea7DK4XD26fKI2Y2lMDiZxBvccyQduhESKg4ajbY
LZk2LwW7dyCQQq3MyEbszgKlpJ8vVgBxn3GIwN5SWd/ZnsBGxSjWYyYf9KLHpc8U361Sbn/UQhAk
kOMd7VMcM2hyFa7t7NJw+ZZ42KfnKsFN+1Lqjhk3acrl/LV87mxk7fIVl3ecL3xiJR9ATeNlr9kH
qB+mJX5I4efacm2YaQ3ZwhPTB23zJGOsvY82cgkX30cieLYfVeD8FSyCYwXAkWwpMq4jUB9UzvaZ
dZ/iPWwHBwRbbplH0yRVXdMO4ha4/gDUa4SIiceyPU+i5XFAvkhAr5VhBxGKj+f8us/RSYkvKXh3
Co5Op7QST/ZZ03rU3y+tvr3mL4O4c3ak2jwPj5LMpsSsMz2sVQGfe0CrxxEF8umwQ0gQebxWQ/8D
yyeubdUmLdhKwdy0Veo123l9NZf3oejOeqcArRPjsHVcdiG+o4lppBmhQjQz8PZHC6bRYfLtVd3G
pfF0cdr0Vv4TFavHiLDMpFuGDnnVHBA3tktH+Y5e2cWW658847Gt/PhC3vi5X1F6cX4GO2INWQ+Z
YonXL5DZFd5JHll+ZafhqBsYLX99zNoNDppj6gOas7klKfB4ouTksoSeC6o2Lu5JwN9xAEw9Lo9r
gklocOjrYO/9djd5LMOOSC/uy578M8eSNfXTl/B868o9DlgJiq++FXqnJ4mA00Q9HU4HHO/qriq+
3MJn/x0SMQyYjgRmO6JXKQzzHUE8RPN0HsQYQ4mGT1nEiIi8OE13JlLZfHNxAp+vgaib98jq6Trv
zzXKkViioThlSi6UvMX49X0RWMRRqNyB6oOv7Ai/SfOTzIurUHC50jv1Y3aUIFqLKLT8jsBx4rVs
UaeqwqVjycdexXf/8HzoaWv7wnu7/scMUDhFDEyQBqQbqsEdTtYerfgQDyUoyT/0YArxBa3oz51U
KuYpyN922z7aCuA7aSH8/DJCSXb+mZjCor9DGHQTXeIJY3GRJtlKUXP5s2b14aOBL4aDHaTGnL0N
13phvfWc7Bp+SFY9b4TtRfw910eh2OnYe2jIH4erU13LlpSKEU5onfg9mgv/5MJjsNQs41h2m372
+JbN4shAYoqN/qfcqK+z6rMCSfxb0IdzKl+Poyzj2I0OI4i4/A8qEfkT9YTi2DMkYONgkM75ehBQ
up4oACbKe+o49CynNoGzvdXdFTdiRWo+qGox5esDgTvJXMS824r+4W9jPuMpEw3y1GbRgPWwgnvp
cMwyGXFfElXriit9FEN0evCXJFZljGjp5Do2/B8edEnDab7SCHfHIXbg+6U6rGp3hixA+yA4fYLA
+BuEmwAWXnny0BmnS/+/HCTDPBtH/vJglK5iorWt2pvSXjW+Y38gc1/l7pVl2dJaPZYgs7rWLNwB
DRNrSXfxg19mPdMd+OT4Da07wEU246yhJIy0alVS5jGfvKCbcmtU7rb5lIqypWH4cEKWrNqcLkVI
1wtJf97TWW+F6VMJlOqomlqPTAKCZozj0T1ygFPZv/cLYOkwIoSqxFkKMmhs0VzuGTPklED1o812
w5YWYMhSN3N/rHh8VSDygWR2mOogb/C+Uj8pf2zi45aZNjitiTUxIBXhp6F+mnsM6NBip+TlcNWd
3YHbEsK1pe3BoE/N23Z1YVwjglOxNdboTe0wVf+vXGXlIojNkG1dBGDlA+Rk/cgBLu7bK8vYoOMw
Qgd3wZjFIP5M1/mIo3+ldB6lCbSnSfln+5RORsnKpO5Zcvb+TV9vaC4ufFZ/8Q1/cu8F9hLHBaC8
imhQO2+EkKgZUMOP/4zBVcZ4v4Q7O44ThIoSzjZI4sbni1fdnbcsFaM2B5UKgWBT9f4MV0r+LsIS
ccVJ2Y5jdnosUHqy39TJRgu2QCPeoyT/gXxYayHiKya7rb7aUE6cBSJjEwWM3hJ2M1nyN2uSNvdZ
2CBq9C7xqBs3yLo2q9IwRrcOQynJWV0E7rWh9VBhYr15HYSfzf552m8dJw6dhtgb+ViwFnKJGRiC
aMY43QMmICUPHhlVc/nmBdIR5E18dc7FIK7sEDlraiqwf3n2oaN8ZncZQlo25X7Td+mYATrFODal
9+juYIseUrwOEIdvHBx3BOiyZL+mYmaHyuQPTdVjlqFHxkqKdKSabWiBWHq6PXTroMvHyIkcUCqQ
kHAp+F908sba8a8XyShUAhy0qTulzHJKD6ygGDPdOw/PZ+exJjtJkbuIVywQRnYteYus9SPqIaFg
xIZVwcMFKfkdw1AVCs2E6RurdhlCcq7khgX/9qTH5AP7l3ZlfeEBGmKVWLbftV+F4HHkqw49tp8c
yk26jLAF90eoQXE1g7SIU0hyV4FKxMfPTsWYhaSrKUQQ89neXMMIMBaLj0Ue+IzfVLIERYRP3Rkx
8aH4IhyrcMQbeu6SeQlcOOpbUvXMrqdhg4OOAYW7RIcM4UWC13HAjPukk0mTFu0IZ4rsqupJw7dw
zm9jem05z7s099eaJbH88I2ewz/eo8rLfUXFKvKRSCaDwcDrJ9XZgHMZOB62etmlQkhMpma00LSj
hZfcyg191uypWAWORt3bvFhXEoP3IOMaQUVGzOFgGgMlWJ3dPiNjnOVO65OX+qW/b3cb7VyLwfpW
TTCGIML203cL/BONYLyFcEAtwWHLa/njgDtyb/KhIMlktUHYxMBW/4j867L997n+PKZYuSvjXjZU
uGtCNkM0zLB8SO1u6xc+iN4OIdYDp9McBZvBGW5W2O3NvUwvwMziB7dRrNlRkm0Xz+5f0kwhuCjo
E8+GtzqyqRa4DxV5xUI4dDJK0y/nBPhed9/Py5bFmKAG7KCk5yR6XjCc+BPGoeK8odu8aPvl/XVZ
jcWX6T1iQgMaEWzS7SlH4HKswIbvhJ+NvxgQwIkFNX2t/AkLczzaxTpjDmH2nFP3rmWxsTTZqery
P99GCI5m3rxCdF/nmYfzpO5L5mz4f61gaqOC0EhILMDaxxSyjAPo+uDZO5LQ2ndp4YJsagEMXbhQ
crCkc5VV0hYg2R/Uv2PxNk/9fHJ3gKiXIYPr6lZIsxy4IUPgu7DLrVRcyr9OoGQ7tZaZyyujIzft
RnFwG0hL6Jd4pfXfxWAYda5aM0MbOHqx5ZAa/09fODijPvjLm9L1PIRS3UsUxp4sa8aGswrgOIoO
rzdJdAHvAPrqpqhzDU3ClOcZJs6SRgzxlL+pEpPD6n/3NzF2UjqJH+qoeiVP6KkyJTFoSf3KCaKC
V812WnEMUTdeu3O+4q8OLwi3wt/ZNCSYGOQ9WeyOzrnZGi49yp+NovOf0EYuQN8Ek1vHo/cWl/04
7VgebZU0RVf9mijocZph2DTtwH/O6pmEEWtnN85aDZkR0/3Xbwui0/2Sls9SKOHdjZY0mcNFtPxz
ZrFcL1IbejP3BpPCJkKPdcKQ9ADrjToS0J1nZa+YyCTDyO57w9J0ZQuEyHG/GFJyQV1NxbSfKuaO
chXlp8gqe1dnB6PiKA0nanP1+68KPHFIG8G74hlRm3aDEmaR0wy4Hj99ZNcdW/MsUrO/jVcDlMq8
7c+cyhKKXB2Ymw7JPy7dft7jDZV7TB4JK4VW5TBd2hG93r5MqvrT4/4my7kVVdPR6PgLDtZnqk9X
lom8DLUM64iI51GjE3oyf3vxSUO52QUwd3Ugklsvt8kUCnzpMJVm9dvFswnBczTdXtr1zsdJJXOk
84XBqqHJU7NbId07mAucLdzM0CEB2NbVSgI6LnS9ho/YkTfgtt/zCvPF/EFLGPYTgyOyXKGtfDGh
lNRBManRxfWRJE9Py0FW6tWICZzoCEMHVVe52YtZFTMt2iPdBVvVsKxY/CI9x4ApL4qNyuGMCTSH
8CwAVBMoxbrJjr8HmgIVGcfeTgDlXtgSmGzTdzbzogDe2+KYdSPeoFg0PgWK1pk17qLyt81p/SDx
a8+M+YZxJvTfre11LKjl6g0w1zTN/G2XeWXW+Te0qa8yubrO0NFDCKAuyfuQJszxZegM/vZDKhLl
7QC13eey2WeP1qW0unr0OB2d3py80AoFMsDQH/5c34XcxPbClSLYhVaRjF862Hv2skiQLoSn5O/j
gMuKke8hQRo1Tn1sq+HzMYlNm7wWhZ+xiPgCkAAL4Sp8ftI94rwl/OSYNeNBUgOnYs/OOtfzBkgb
ThTbQ/XggisFFvGXz3lRJTKfJ0XEpwWP/3hHmhl81URew+BIDh0pmrWSxrTM29jRaCkY7lF6oNM4
eG0v7FN/igfh8wEtz6tUO/B8ip8vF/to2hqS6E7Wi4ONVBL1VO6PdjowGDp6Wxz32ySbCLqIndog
okeezUKAMZNXxkfo8Pb3Q/KHft5Gw6dXJnVYkmmUuHjSOJUG3/vLlxs1PJS6vMMvwdceaY0k3DcT
2IoSIbOQRvLLscePzOBNoIdzmillf9OrqKN9QPkilNZHWBWhqXsFKvHS+lBDl8ESfYFd4nPg2gI3
39LyRC+HQv45YeukUmG3v0lXaYAd7c39r+YT0QacAREJenGBYfIGkoY+0sOx25rXXDbm/IgnHkG8
+CeWH4Tdi92svruVi5wQCLvZOUUTj0Bfi1X541ZCwJD40W1s3ZMBYsuQ5afgoP7MALQN6vce/pTG
fniQ8JgIG50kZuOPIhOE6gAgT6bC4r5wcf9GTzOZCWweAcoICdoq/k0f5TTB2Ok+kVL86lWnA75d
aQfCpoapPJdrCaYrblKP7xwLugXDuVVqe32mnQ7q4GsrHLYIQq0Q0fZrjQsF6FQTUgJHXh7MMYOY
cbNreoSyC7KPcLFraK99BVe/DQpTVsUb44bEf9u0CdxN1yluvjEc63Xtjq0QQgz01hyz6HyBwdYr
vl6yfVArm4XK5bF+FuWWQH/tNXWqXeULupQgOSmZ9tQuRghMyD95n5TeJyNnM8dOZDMJ63BQLSpe
lue1BlqWjEA4/kPtOuMFtxHXSEOfsU4FGJ3ryoQZoD21vvL1gP7X4WBzZ14YQRNhwdENICqMauSs
UoBqzG0ga8hdVi+k2ncH1dJiwIj+lJd2plvxQYXcmEeWg0vzyaqQjTNEms7tguUf3r6x1J30bsIE
kn+Zc/MENvr39FQpwke0Qb7kjfP/j8H+PGvb5XmRpFM7dWHwHSEHFffdv25IVdVWw+eFNuHNyZ7o
LJljP4YZ9hbcTYxZBeKUtJUqyAaXqIhj0P+4KSqkNDzDXJSyETt5sRBuNc/rTkUERNJJQeBuE4Is
TIwjfPsSetECJXrTxTL/MgtFiE8RCjzigvHXlCwH7OHRs9U3TIJ+8FdTsxKgsc0TBmQaINFNBObo
XP7dMchBp2+To4c5WKQoQt+cPMGGCS8Pe+R97RwUkoIIM6iaDH3vcbSBIrlmBuEX5HBBIVmBrNuy
EZe8lsMpKhJ3a6DnGSSKKcgehD/dGC640NzUagCf45GH84r9+hIN/nrKIJ6lSW5WbUgeJ5eaWiME
dJBDUr9jHYWPQIZl4p4+KZw9UfdtMUozDbBp8LXv/SZnsROUGS7JmjUnxYm5KzNlwyLVyOrfCRdh
T8b55f8LKwwnMzM73f6WyEwE6PjLkjoDzbZ0LeemnksLedpkbSnbSZObLNiT9UKTr9DAZi0yJTpL
ldIn2K3Cbs7uMZj+asc2eKzwyZXPksv+VY02TR/ByE2p3sub106pV1zLYV2i4hmG0KDQGu6ILbnr
qLyEwqRcmkQasTSWOi3LwNTmS8mb2NZrQ+5RsLuGpcM+j3YRah7wrNv/JaLrGqMZIZb9rcFuAfj9
+9RMmpOT/Cy8B1ddVS1yEL21aGEbJ2vcRx4o/2WtwLkNFlq7Agcf+pEiXtedoCdfOQfmBWj6U3q1
4vtVLLM54USmf0NXb9hQc4PsKnMdXhhjIHkwczcqeBFnWKJch+eWxneTc8PfEqjGcB+00FL6oxqa
/aNONNRwEOL+e/G2evVZ0Y5mnFX09MW9lIb2f+fUboNZQckU+fLQhUtQgv0yYo/0YCUYTv1neXBk
fy/3yqYqKU8r3fnbscOSdjm9F81Ib8HYpiMl9Zc7EzCIuCpCW5hbvG827TPvxnxSmHadx2z/1hxS
3Flb77kQbXQZAmlFBcxQI+blxYUe8CWmCFF5vL+V9Qtpn/f940hojk5keCtvFGuzgMixPlq6hlaq
mxyU1P0eypiFXaTi714eh3wuyL78kvfhWZZx32CWEKlleh90pI6TZOw4rB6J88lBZu24wIIsVEO6
tuFHEos/QJxtYk3fPqypwDQCQUyQ9viTHNXRQ99csKrBJUNVpLY0pGFzwxn6slp5j9QGIWdDngNE
gXBnMdlmd9AcsqyoEFR3K5HVB9lKnKFT4yJAjYFGlmieuwlDZDcek+eQtJeoZo0E567XbLdtl8HP
o1Dx1Mzws0JS8spPIi2PqVlPd4WXNh1i4LOjpffIMLv/bUEjaA5CrBziPnQH/WXZ5U8Lp1cDqPvm
IAN9h6iXci9NrSC/pdkOrQSjoejknTG3itNzsqYDmh5tMPVOlxvcvQQU55su0RGiTX+A3JGdgaUS
/8G7kyot6sbiqQKkgyYJEh4wejH1z5rE78YdJ3fhMa9SJoinG/8FTUWrlwtonlm1CdlHs00IafCk
IDC3XsVPwCAFIEKRFc4C87OjFx4/EoT/pQ0x4jdezarhetV1566NRs8L1UPqtRGytSANaWycQ8Y3
Y/dqM1Lgn+LjuyNxLKD2lJrsA5RP2WieZu4SEuTCdYjc97S4Iw3mTc1FBNxTAMFyzj1+LRO3E34M
z05xri5aB9SVzI5ubN3vyQd+y/swpoqCzS3pInQY3+W+ND2/gtlRS6GT0Ttwqv8QjdPH9v2vrPFl
DPX/RnN7zp5xEYmsZX6YJxKg/v11cCRUa/0TUtMA0VyZMcSu1vZF6g4W9VLQ45bCPE7vzEBVYd7Y
OpnLvlqYqIuruse3KVaXBlWDQWLnuL75iGmHzCelAz4rXsBRDVKssZC+V2EAFPDLCWU1wp1MsoWx
UAirgwgg7ENDi0Zzvc6GsPBegIPykj2HSYFnPFwMOacz6wrksWsz5rrrhnNeDJKUJA9GGzLjUuxq
FIiv6Ju0WUskeFlbiniZK4KjYPkJF0S/kT/KKz5vDs8V9ftZTj0Y6U2l8slHXDp+agKqzxAqDqiC
wGnD23Bv8baqcj8C1J2r+I1sppnZXDYrucWKm1G8XsIX4vHIUERtJXpXlc4Lk+dk0ouiM5BypzZD
C+50WOc5yUJ3dxh+MBcc7kY4ALzfy7EtEJ2WKwwIOH942x5xmCXNO0DRXFd2xm8LB1qSuYB0pOuA
N8ZfJevN3EpO1mkSda9P+kb2W/fYNOlUmq2hphLOcAuf2YGWm21KDY9fs+5lIgJVvc8tO85UZZzj
qFpHc0/LEnEALUyHii4FYrhfo9IuQ72BFxEG54uNj0q12afML1Ax9rFOUYUZe0MSTjy6UhXzzLu9
G10FtOugl+B1aD0W9ga/9jXKVE/ODdaYx/Vm1JKbO7ZEEmrXuorQ2QENe8lQMRbxPIYu4eq1wy32
fRO8JfAxYnqZ1xEMYjLxpvfvHC4RKmnSOBSyd8KBS+YVx/gYZ12xKUv9UxVYlH/CZE3YwV6OPKud
E29xlVEQcBKjfGZLvpFZ18u0As8lCV71uBocjjIJX46YLLNVH8kTNXU5+RQ5vwgaBqQODwoxuQm2
w+z21Y9wpXv4GjbOqt3xDWBeuBcUDmtVvz6NR91145WlHaDuINkjVMQ0+hB0+pVxx0IloZTZBZXG
IepON5cGAAdyKuj9RWNXOFMEwQ/wIEwUpKJsHCQYEmoFBTXGo4stKrOPR5tm2xwvnQB4jHicHqW2
oQ2jiqC9WUyl5WSlflQmIKXhTV8KbnqiH0s4cNg6ho/jhsEXxwWZUC+b7CWwZQ/UDjqbWZQsQW1J
YC/nklk+JU4Dm6w0+dSsqWWiQVhp99Ldh8ZgINxqfsVMbPwf9Zktks+rqBxdE/RJeOWwYTAN0rYj
D2yF+NdRlg5/HIq34pdYL+SxLlGqrNC897unNopqb3E9JCih01V8U3Ng/RY6qLG2bB1/BHUA4qwR
8GoHEBInruHGH0wixvOyFcRPxTLdoCz8DLNm8UzWOpwYfxBHpvEFNt1hDkXORqXPA6Q1fed1wQXY
YKWvj+3qAVQGzSk4QCXNi36jjgdbAqqyiFr/peH3StMh2gJMyZqVIdltyO6sZG4CNgzYxQ6hBPk6
ibMi/rGn6OgRwqBoy/h76Ser68xOMi7UvHXRT1/3Uho6Qt6CSvBihFshtKY8Me5HuolNEUrQt+gK
JBJfYtUAAbMifq7LIKxum+O5iCNyxw6JPIj/VJSB9R3/+mQyLZrA1Ac+lPm+31n8HkoKK7/uqvte
lszdTjXboItmDRIOomYkXD3GxPYX7GHFG/uN8saPNio1gBEvaK0q1hq6Td5tNuv1X/99hThhA9qi
Z8uEEsd/uzEJWVN81I2WrxhpBjTw9xzV1eT7VUTnbdjqtPxqvdH/QtzYWSCgR/xwXL7HxW4pMdE7
+FVK/CKfLVpf/PzNuwXsbN34yxjYqBfEZWe2Is3pAt6tD9sda3lWnohWU9fqxxz6lc8jkgSIl3LN
+bofzVdPyiTQLvakC6xwoNrDQRJtQqIbE9BJTcrbjidfCljkr6EJfhmHHBrLcVxObUH+T+fClFc4
FrA/tQfkSzlQXpHIGhLv+eCDesgdcoXIIF3YDim5XRqm2UFb+4tbXDKhfVwV/i6jX2a/CPzdROCE
Fi523mf1mwQFtwIMc5iyQmdYtmtgPZGE9B6cTmWi8kpJEOaTyX7dD3XOW8yEQFtJoR9vJWyyT54Y
CwQyc5tTjLbql78shq3jg78Yj43HccCEVeMOJKnzNmzbEHXDi+csibDUiCKvaNR+yWs/Q8YNE3KZ
C+OOfzR6oC/IlfFIf4O+sULnXNZUsw3zZSvCOkcuMxGp0HaB3XE8j9ecSlrNfaMz5v49LmFL8nDO
sfb+GA5Tr9gorLQ5B2kMtvVYOh/OXwLtCEst0EANtOb7fQ70BcYiST/i5wpw6Vnmi4zR268064yM
+EwWHpLvkVAzHomL0nU3JSH1KMCc+SIJOK5IY7RzsayxL7RTpLHJieGy+Q5amNAjtfdTPRBulyJ3
U6/UoQLMWDI3lXPOBtEV26S8hIiN2inUIFOPBY8qKFVCFDsw6O6DbbXl7tiQMMcyM43s9lThJcxx
GhtLvDOfhFU9IjMh1XRyEW9znJj5r+NRtevM5q/wlmtIJ53ylfHmdZ3TKermKB5dHzLSyZ8Qu9hx
FWs1KXtWJ84jZg6+RqyHdMFAs/DPRyODE9KVesmIlpq3vFE+KhGXIAbX+xaszpQ7ws+htWI11t+n
P/VryuAA8R+YnODMrHFKDM1uEoWm5plzppWCmD+bBqMSLmJNxuQwR1jbqTzmZKWX5V2gcY9Vek39
D9bTSPNyLH3GbORiRrtMOV9/+vpnPGxT5RJ0UB4sZaw16KCViiauIGVAk5nZ3fIhNf6JPs2TNMLL
9lLzrO7PKClNDwnwUC2qWFBXF/VG6VDJ51eGdNDAeF6GK1oIE28V+LC08b2qtXwtpYUnthMxaZEJ
bx8qTXQxKM8j8PNSpy/P0q4mYLj9JQCY7m4k295jzmXfZEwv0kUvRAFToCst+TChTZQo31KhC82a
tAtshwzgsFADHzM3ELRiBPgJk7xx9gWW7+ZtipFcyG1yBP5CsGpJC15yrtbdQ6feKqEqLtI8HQWR
EwX/NhQZfP8FPNRCv8x0boigL7ZHn0NbHLzJqOnuxuHdtPfzsc3YItH9VRQR/JUVezxL45gm8KVD
QCGZ0w1Y1PFEKGwXewe8W4vAd1Kdbf+wanR7jwLWJQc54vnR5q37/7bz2dfQ9YuyZx71Xhxh5IK9
/wqIGa4SD2ENhOOQ6XQx8w2+W0jkZImZQpbOmnufFNIHejWErMoIiP4yP2APMZj3K8shSJgDw1OX
C6JXbZfG/U/ZsyQEGiblNQye+Ig9VwX6PYTx8Q6z+dh3md/7SMMZ/jPBvTIAEfFumAv9G8laI4n/
YoRCZ+AzO8sAOl2JL2tfB5pIzqsttm+hI1OhhxcmDl21nOlwkJOtpW74lW66RhGCh7ABTo/MQj+c
Shbfgov7jNr/Uwrkp2zIN29wnGPHCIpBfp3yjQIo/nByxrKtOMwNe+UBspgIsDUM2HfgkA4rqLjw
HmffHkzTLnSO21HS5H427hgvEim1G7DOgOfgUxwHerzytzVfUXh3tFMRc+v4UQ9cddT5FJuoS0Gf
7BIknSzXT9XehPgqs/yAhd2pBueH/JD/eI9W0PUM3TvPLHFuukHAvZeot0ThAl839xDbS9nEMQq/
yt/0ghOCsypsh9DNxg8JK2E+AR2FUH2am72kCJQM7XXKZZqt4GUwFFPyM/xXgnU2mACMya4BQV2T
Qbr+nqKmuoFjL6vB+gMNhmCrTJB4tT1PauIuajfSLmY814Z5rSXwlXPJTIc1gogy065fuvFvjDI1
GuobzcuNX9Otjz3/32k8S78JJfJp+k9D40BCVgHRdmBiBCpYb+f/j1s0NIkWzg1DbMv/HesUjGGW
1gxJHpnfrs1puAKWBzEQ31Itc0jxvWgTkV/cn/B7owVqSdY9blvSeGfWPW652cNfRdXaG6pa7peO
yoEg1WmSAFN+4GY6RMXjEWixS6f9Y8BX8Ns7xWh/Jb59oluPWmCJ1blp4shc2nQ5va4L3rGxjC3g
X8TidtmAMkAQfbAfT3Upc7UQoTmn6JZOpqK984J7i2krZEBXJvjaNiKGZSz4lGKaNtI3y6xr+9gs
EqM9Cw7yZuIn2xdz9x3Al5Id532k+iNq0rNyqP95v/7mdxB3NPXVtSSQnINpVg1Giog1ln5XVWBk
g6+W2yMwsSxrfsDNOjgDt76/JH99C6CjYJPV++FfTM7s8Wnf4x78fs0yCya+u5Lnp1y3g9UEGHUl
K9B3+tx2BimX4+h1sLva4ssWYafl5AYxjldyONx/PxAM1S2oNdSW7O+mSF2uLMkwBHFGdFLaM+cp
2XoNxtk00Y5XrWGK/NgkRi0DjhbI07F49xMBlx+nPqxqJj2hst2AGn89KRFqF8oKCK0LA4IR+UE+
iAdgaTVBC96/+mRdmwUGqvOOrjfm5oHHpbc5nv3jhl6U2WPt6HUsKmuKRsov8tu4WfFeMYgPIdjo
eTj54NO7iN/e7tO2VVWD+SsNGO2e25opb+XdyFVPcKDL9WI7cQoDZdtkVyEVC0XJnqOADCsPjypd
UiZuPedRmq2/3f9liI0DSQ8IFBfscFo0RxYSJYcUvDxYRi2QkH5fl/bAaQe1TuAbmqomqG6GD0Ie
eXUPuWqd1dFXO1WjejpX5qW4SNXQqHrV5bJS/4/2+SAYgjkpR3MCJg+jCon0P+jNExrazn6hI/S6
emb8YCxn4mY+YwNu6JQuRvKwo02aWTUNKsnoj4OYz89B86rHJVKkyiNwh1GhIzl8GOxhAeVsJMpK
iyn9M7dRRzUryFewKw/ZcPCNQR/OjPTdCzUYTDvT9SBICoWuNfARIB200/1JGpoMsHnnR5Z4nYwR
Mh0cWjShjQxyXemCPhF+uwVWCfl+JN9JitKgohj1sM5xfwVFop7mLeUWroUk9nnbqR1OHGG+n15v
AjbRq1PQiB89PEVQG0Y2PfZhNlv4USs4exFz4ZsDcNBf47xehqk57h2YWxPLhHS5nQwR58Q7dmRb
+bNRhbA8K2QOEdIRwTxvUaNzD4YK2nK/hptGwAVE4fYii/FpgLE68h/JRuMWpmuOxKbLgGDKXhQ2
ErhOfmGF2zLABpgBQbMNBvaQ7l1HsD8uvhXybyemYOOrpu7hT3w0tSmFubyw/Tg8BuBuaMhjSYcE
pkAWiybDPIszv8kLXZg1m6PRGIK8V4aWC/L6NsuLMNJY2ZjyGNN5wMfZpytfhkL6qMEyYNw1khid
cNT72gEMm1LTpybq/0CMbOYrvjCaDOQTLkvBPVx43mYBHhzHnwzDd/dq5G/XZ2MpD7qDehhbP3vj
iE1pb95CdB0ydjEMzDmyNEztLfDIyN/mFHIYw51dSPFnWPJU33Sxlck9ni7T+dgaWDUV7EHjYHCu
pAKgFJ4KaMiE6KXJpVVV1p2f0hO6IlWv35jgCK7ksVlyXzIES0+5uEYdqUGZNYAIccvE3bmW/nVm
GeV0w2P3cit+vIpDi0n8+KiXDz5w1Fw6ilAcmwOvyBGASAv9qewBqJ6exNKfe01E4WxeXpCYgpyA
YppqpxSXqDfo80BQ1eUUuHwNQLiEdnA/+WFnPAiFAWoRtOFLvZjH7yopxq3gv4tjI+mPo1a/HFHY
AAuE5I/run/0Nh166/QUw+pDOtoHNE+nZGtqR4dAlE/03WJZfvVO+HE0EdIvV5S/18guSarYXYi5
Xc8JjJ7E966SwOnxMF/DZubGqiJWtG1zEvvo4ab1cn7nW3tPRpaXvyoW6y78qQrvqAvZDa3/SETb
/nMQQtkesGdmwPJTGLN1FZkEniTnvnt+GpIFsSAYGT4LaUki/zJ8uxDLqJA5daFZC5wmmck6PsS8
zx1N2tWI0d+Bbm9kJQ+6QXaPIKxH3RGB8WsnCw2gHhdE3iVw/a0zexpydXbDRRIou/eOkBrjIgi5
dqsdkFeMLc4KKqmADlCA5BwN2RL9WiAooaBYWXzQOTRy9YvMIG5O4YstrsniWbxa3Ukgiic5Z66L
Qw+HSscF5A5tOOjRSmjPnoTfoe40D0Lav1JGiS7+LhV7JR9D7nA9nb57xDase4W61dFDMWN6++sT
Q6T3yv8yIAxxIbqzafQ9Jw++W7p4PvlWfJl6tCnR3qTQAOADEyLuTMGGaYEwdT2O5VZJk0f2iSm7
g9g3lSbreGzKva133Wb7A/25ODJw4aPpPhqCau/Y118eUizH45hbTu+jZF3r+RSyHJ613TgidCpI
iX0xeLz3637rcLV666fHbb8BvScLEjF0puZuNnh/sEuWc4MGLXQf1Fql2WgJknykuBFTgGXrU+jk
kDAMyw73UHK7T8GdHDPUtHEF8CuIEBTVyfJyP5oWm0oYeIcL7smIwoGLYaneDi/d9zgMnsk5gx+p
XgktYxRdmonTjg2VmYV9cCLTdZ8XKSmH6g9h40iQAQ3DQ2wnpyR5QH1z39pXlOdt4blR7p+YxXIB
KSq/rZVpMTvSbKPcRIUAeY4oV31kj8E5NFg7huJQS8p7E3DAIKNvmpqDoj6Ki8R2/OEW8BcLqmGD
0EtC8uogY6lLzvFFnLSzrg+fY546tiggBtnR1J1SR8xt6hYlA0UTE77V0H1bzGzM7ocIsvesPblx
4j1KGmLnkCcoX/cu1cJGTtjLXf8RTSpM/IPLnr75wjzR5Abwq1EXFdYfglLXifBBW+kDCYHlzjTQ
V+pcD2M1odpY7Ji24ASa8Uk8GlD6nXaWGyOGC8FDNpeX24hgy4Ae/r4fKqY2/bQ8gZO/QlEQQ9dF
Ni9e97GJBX5i0aFmjuOO2hz/yV3T97aG8TT05hlUg2kbWZhMpnq5fi7LaxuamdlcXah0qaNF3/w8
dAVP5JdfKFX/yd9Kt813knp+Cv0OpB4XAN+XkN1TpCk+W/FYhbcY3/sVEFF23Czhuy2ezaub6dmH
QknAH6WtCO8wqkx9lj85MopS5MGbHGKATtFXixwdRaTJpg5sOToZ+89brCgcwvHooVEckV+dafQT
7Z4fnB5v9L25FwbmDs0wMTPkYXEVdpURGg5NNk0ybqm1xGenv4enuMA8++Zs/96QL51kIRfGba9r
7XM5abIUhdLPmEMP5h4sW737vH7k2DRm63oVW9158SrPcZGAiHXWGLblMs/9VW/x3b3CJX1xOPkI
u9EO7gx8LxXFFlHuZZcamSPNdtPG0IIt5H3zwjQVMDT6DmfX5cryrwG9p7m/QnIXc1T5r2OWRb3a
9IiuycXgs9tI/u1m6GXWdVj/u73s9J83WVaRGDR0ABgWj3m4Hz4Ndj2/IjtMERamS7HaEoQNk12P
woDzT6GMwcWhcW9C7J6Uc6cC2SFPzqA2zuUfU+VgyhsAl1fUIBb5zKH3RPhhTPiwU3v2ylP+9CTg
7IzML3EqA4Re/avkTUF/8ol1n3L5ySMGf9YAhEOIxBc60ExCUUxn9giJACmrgJR1oNWMnhNyuksv
w8JK4PtddrTv3UYT4ZQSvZ3uxAToNNGZJKl5UStCLonUEMOgkeCFbyOY9gpTkp008X084ZEBw8Bj
8jDAJl3kr5tHmj65Y69/7fzxdCwIfDeiGpTd4xCG+tYG19MXCbvDZlNAnkvP2faYEnc8yA2jSoif
7OFVBcLbtIIQTRiBg4DQXwIVAUcDrXodF39oFJGIGvF0Izvsh/Sjc3XDTOYYw41qSb9lBrf54sOv
9AUP5UAxpJlUwmY0zrx7cUInlJSso8quhlrm/4iNr8r7YejsuiP2Ht/oN9w09yovFEAU5SgAQrDF
EXpEJtCwfrJrvd3ph2VHAAfVBBKCsofClXix4zGCXnekXcZgEvrNqD9qzVUHsrTWsm0XPjlt/uz+
pIeQ5NyXp4Ysoo2VA8+MR8bFcPePA3+bNSeaVU+cor5bwLRrtkLJfhc6CSQAKnjjy5B3PKJC171Z
dh10WpLegPZMaeIW7UW7Sp7XBvZmWA/5A3bbSA2C9JQOJw5uMnLZfiwuIDDTNIBDjhTYvry8bs19
U4qdDZfWG0I5xD3FGRYrYy2L6tYIXanBLB0=
`protect end_protected
