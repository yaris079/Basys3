`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qPR32iAhVW5nP/IUjtwdRLQBtgJqxJzSqoiDIPLucIDFmICtc8aML/E9sKf2tBrTwPkHo/I+shdH
msjV/NIPQg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Tr0uQSwQroNXEILaQTSdNA9EgS/bDuzi7aPBEC9G78fNFiu2YsUXpZg0tNiC1/vmKumJ6rtG/Jm2
DJq9jCDrNgYLzmWSdaU2ptLfB6H70Ntn4uuUzW2GF3tHVu3erdyWcfpklN/i/Nx4LlBWWgorqtc8
S3Eb2RfF3nuTT9KMWpo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F6VtPK9AjXMao2TUJbWUTOGLjDqdj/GF6SnZumVLXPOzta5XzJlcf52Lc5xp68Tyi+uc+Nk6B768
3SM0xqVXBnTfhWi4AtBfeOmjB8bfgoFjeu2sJ1GXfbLQGDq+g5eMJN5iqpJFOFShm950qKi/mFhz
Ovx8qBZgTYvRJx6Blx0qRQ7Hld9HdPWchZUAPFIW++zC1DVbQ8t849seWiMCFYPPapSqB0UsnzXy
XsFmn5mtHPW1RX6TysWYB3EFv7dZYt0cOORr6LP39nmD+p0ABk5L4HAPHGQS0y1SzO7RBc5M8qMH
Y+7nUAmfT+6i5J7vBLOkFfE9BLcfnAAdwQExXw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
doenq8fkJWKFJyBcxK8QYNDIfLIzfPVmQWmgEojLwd9ippXxeZ3jNeVWFP+pO9/96Y2ZQIgVNvyV
titW0Ixw6cxXtovvHuh6BZoohDhkQkULesFOG1ctmP60NOJQR2DfdpAP9HBvlkGsq2UMvQTeNzO8
+2XPD4CtbUmaZGB4Zz0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
edeV6x8zqofGotof6FwQEUU4byYtz7HsGiaOpzNUeD3JACRWYPaUFc7o/OVDhHEID0biJkby4Qiz
rN/vTyExoECYAMSu6A+fT+I9ehYaW9YPybYysiWZsuOdhTSLrzFTkRDJlNWtEpCHXDAxlN3GwjsM
50UU4W/FNSoO2w9A/JNd5EpS0hs9pELbEnjNC+AZIY6t7MFDPKOifhtGFfMtTIegu+xbwlsgF5KC
ztpymepgw/45Ky4tvg9V4SGhUvJoMJEcrJlMn5YycwLmPIk2Uvmgo2IVQRSJCD7vr61KFJYqAeil
UeomP0AvtzkuOK1lyNKuMHOiLL1tF8/aWM/4mA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22592)
`protect data_block
w04VKlqe5v8x3GOHaePDBE6mQv2JAKXw6hrv1pCK+1XPvbpluw6qJDNdBcvlRZv/2Rp9+wnlQUN3
/NL79FQYhBHQ29tACELsn4p3rsi6Ho+1lUqO78HkZAGKnd5CU943RZSQTFP7vtBUhhKpQ90Px0lg
L++RhCDgptzGWAeLQwGn8RzYDwMMewA86Qd1v5iK2cXo42Eela3kZOtSNf3AnjfG2Vg+FCbf5OBK
BTQK8xottyGF8mkOSvZh7Fxwt6TGxHE7c+asUbxF1/QvLrwZVbvWTQCMh3y3dZZt5Ij9YquN1j3X
/mrVmnSDk5OCPIOavRk/eV7tbdrX4AMAUxtKuFOe0BFBumFhCMi4V3AoV13YNwvKse71EvR5vVMM
nGkCp8+Yp1bhMv+agTbpgUyZixmsOZDSsX9kpj2V20dHGaW7SKugI4NXGjBGQRmujDVRJWpdy1vx
HwPfdNEan5/1ZW6CIoKJn0SH5GRjLEqouLOZLxTHj6uTdiHOZpzIHiTB0OKI5N5MDMRNm92sEnht
beBlqE7s8anUPX61dTvbcBsiVSSWmX/sIOcITAy+bXmae6jagLYho69Yw8d9cTQ9FfT+R/GA/9yN
sMKc0RDbvNgrH0uABUCqXoudxHupWFNQi4WpN/XDF8zLXBH0Wydb4ZWlnxRqlobS01BV5UDgIarX
LoDvAF6tK8RaS1/Gr939kwrZ5ICKCSElWTaGxNVxxIuREJKq9zPb1ROnW5UMY2PQUaOFeVMYXU0P
TYVZGhw7wscxulfApfsZTZjF1vf1kNOoLInwgtmgBsU7CelMSp4yRJnBXhAKhPpUq24Z4kQftSL5
YcqU5PLYiFiWN63+6aqCsClpX/leHkvsH+G3E6rL6+V5HzLh1f0q+wBSKL6T0BGbqqqC7KKY1gCz
Gbj6bBzZFG7kD8p1tTKaHiVL0GVfGgeuJAhSyIeQZnKYgGTlwm5gtZJAqyEbDQiCNs6bTAlpoUoX
5ZEwkqq6VX/k3d7xxCzx7meExd2vI/j441ilaGfdQtrCNqtLi6Clwi8f0sdpswEOp0eCFQSNK7ct
EohV30qv8mBfDMDdoQZSrX6VgQ2QFR4fVa9exWT1NTOmh93h0sHuKSRpSW7Y4QijP0SER+kBkjJU
KML9TY0Ju0uEaSFlNjfAtYx2e44oioSLb9zfBi0UIl6wnJwUe6Pidh8tT6SUW1EBaF2U4JQ7+Vj9
M8zhi6/MQfu4Ox3NL4Z+EnikCBpI3R50SE64Efd/4NjespiQ9dPWZdRwsN5zVsk12ykSW52q382K
P+fUdPOgPHeygWuWVPt3c9KVJWHLjT/481O3hKkXQjkz1ZLLe+JfFj+q+R4i/IxTqOXz6LYarcam
fA2KS8L5Gk2l5LxF7TPAdP8thKwr8ZuP6hMRBRqB4AyCocfIDFRNbnZ7oirUWlhkwnshgFVA0lt/
prwPHKdxY5Fdycfb6MHVWJ2VmIK7P5I4WNLQ8aU3kHevhPEi/uYcfiZxEMJoj8TfYezuS922GQ6J
nFsdgIxw5wV+wx+jPxBNu1qXBIH/gVtdvA3LYUPZRDwXv2vDcdUtnWTtnMZPQC/CpTbRaXunAl5O
mQqeBix24ONG4Svj9qghpTfvqFvt/CLNdg41Y31k3l0OC0BjL7EKpgqitpjUy5CqS2b7vKM77zAq
/uFBCbE8HWRpPktj7bOW2IHmk5ahM4p0n3xM5RH3XLgtIDT45a7HuZIHPE4rofa8qA/Fzwl+JEA9
iNYBtzpXKABSDILci2sx0RjxXUA3qo589HplW5EMjJb49m9mkoyJTs1tUbZ6BL/snXqRQynwKIqO
R+5jpxYw95Km9OjKaai2p/098ZM6oz1TVKOAckR4Y4QlzNJM+qXHIkM8kVn8ltwGMmMrDXvkhZUw
iGZJkwpiw/livbMrICST+n3zLSMsA18TBdXDteRFnC6Td3KqLV7TxjH9nne0SiaximImZWUUFkb4
uUegL5+Ag70IPjhiAC817cBgzCZio1ykHad3A408Ew0gU7OLCvJ5nBzA9zEMu9QGR24nQOUDcRU5
zdUiQAWxnrFZtf3HsNiuMEHUGgRkzE3wNa5qDM9ER0pBLI+iw49weFC9oRtooc/EzpvOdhGr5L9U
ml3qxr2dCb8yN3EqN+977/FC5mbgkdqRHN53mClSNUO0WvZv/juCj4Rw/RcOZnTlhz/f7oVUx9Vq
Lshyq8iW6o6OSHE5SuBzunoTEogUUasGh7HrPqUJ0vdHyLWUMK0FJ8H+p8y38bBetUCiQg4J04P8
qTjV1kh8cm1gZYS3aOpT9Tiu0mSJgnDqMsizIrXMvdzJPXQVFz+CctsOdPkIrAAMsz56Mc6SYitU
aBKOZYUmfqZS4wdGhkw6sJ4RlCvJSBiH+2UquMot8rI6PeAMJdeerwL2y+2oNs62ii4PKj7+MjHR
uD/mp4E3XSEq+lJs30CyfU/MlFG4CTxUf3k21kAs7UW6XvY0VpFI7ShlFUq3s6qfJEldkbtUZZEX
gxu2PrbrqygeknQnS90azzDTRNysuDZTyZJHa0DiTqw4nSB3L0mfLoeWET9i+058vzh+Z2ICtzk+
LFcfT2EGleZk4k5L1K0Xi6bT/oN3EgaWCbPD/fh1oZ6S8S0M+sCgt6qq77iFk5hMaMGICOAF1aFU
FJYaNyOCoY31tnzuraunjbcP9+r8fF4MMKbAAXRd0Tg0Zz5hzwW5/xrLexisGxLCq4qvUzA0g2My
+mW7z/8kN7HBfDn6C884Us1EiX4q63jKYtlWN17eP7Gn3PGbkV9NHPuBkPP/lYMp4qGTieC6zUWp
1ce+BiJAXSkO6L+Hd5hyqcT395vNQfD1uIZFwaiGu7gqFLT8vzpiBo7G7LWOdnz3WvlLLHgdNnwi
Go7u5+c7Q0IlG+VMmAm/UWIgu0Yq63NroAXG7gMba0KNXLVDeX+olirYsivM/kj6y8BQmEOP/jfA
T4MyfwGlfnwc1ImKbhTS51Aaurut9eSDcJxGr9CfiAkfI7U4vmeY9K9aVv0ledGdrPMvudajCumm
L/o9bzFjuF/SgdL1VwnJeAjd7yG6Tw7I9pR8iwnwbUh/rNZ4h86dqt8p4/bnpaTj0drHUJQ4rdt3
AaZZBunaNODziu9j7mbYNzZHpCKHLKJksMvnTgZMianm4z23t3LuOcrS8a9L+G1LOrd0ohVZEBFo
/8rjPdgH4X0YLRnqLClqTaadgkN+cLsqPlD0GpjRvzFRGuvIMBkCqC/vIB0b3msdpxxF/EG0SA/w
cttr/1j42ENIMDbn3M6z1RPD1E1qxFa4Af7HxDzv41jkzOZMMjdt0rXz5/Z8YUY6USfb8GsEA6PG
O6J9V0LvjofGDl9dqn06CxcEGmLwozAKh9DwZs19J0gkpcVpxGaYbyat5V/mWF5iVU0V0AKV9jMV
U/1TwTWXOAqcog4d73SRpq8IbuWHZGc05TLgO1aNlD4wndRM470wMv+et6GYcHsL5+QBJuwI00wQ
Oaa/nXtbpNhaa3U/ZXi9smxgYPHGoNw0S9gXj25lEe6rVWT02w50UjYu/fXr2f8WN/tWmQpOJ+Ax
grrlNRYxeKXOnSshuu+t1OEObhCY4uf61j4QTEMHC1FTEw1n0dCpBCmbLQI+SIxpfphkDVzXH2cV
4ZGUl62lUfMKvjjXBdsoOd4NNAoMDx5/oKFPs1LFdSJG0eQZCaYhp4bHvkp0I9MzfKBJwYLlIWmo
d90eayHwKuWZmepBP6SVx/178ofk8v7dPxoIiO+fcWECYyMGxxlA4YZownTDtObiV+RLYuIr6swg
fV4zc/GhsvrxKXfmg//XeusVZqkUGqQR95K7Sl1NE59jBuP8kq5lqXoeZ5RT0VlgVKMidWBHs+Ps
G9rpJ7sIKcvC0tRdQjBKRIKZXB1qkmt7B/+SFVXXy0j9G54Oe5+/QcTRl0exS8eM8KHaHxmjjMmM
hF8a6efWcPzDKcoN23Z29HkJ1QR3rreliV02kSfLb0CPHAYmZnK8aRISfgoZvM9HNrFO+wHURMPJ
rGH/9+9ShrsHe+6eukvEPyERR6BJIoXpNHlxDALOf9tPfuJMSkTQ+dF94Z2LDgJe0vuvMRtWzH1t
CUWyPWjwGyxo8CqxH9773JuuJ2OKZDUFEUuVtqFEnteEjT8n6EEdYN726pNycGWRlosqehdUvmVi
8ZDtE1M54B0dvXVOFlrf4ZQSfxk9CvI5ASXGKnaKt+wUSZzZRANvQ26j8SlRrWrZwfKU7a/Z3Ewn
cTOhFOdtDODXVX7xPxB+cyRkMNfYVgYyXZr6+ncx5SGFHDcr0mJ/rZwKCNkGk4KJUu1JNfDbXAue
EebjaIu+eZ1Ul07QvLQW4tK7b9DjDyiLJ9zRvaiXkmeY3CyhMpYoTzpjvEKAeYnBlG4feG7MJQYl
ogrnj5HM7DBVLLYGa1Lw5UTvfQfreBmC6mwH4cJJPvhIYhmIhZzaCC6cxxvN9QEFl6MmTt5aXDFJ
Xn91tAZO0O0nQY+4/BzNKdfOyhK5si8XXZcV019EzygyU2n/FBuMnftgcjnW8mO7Bsj/vZ4UFpJR
PjNGHkpw1OTY5jg5vLdb/PvkH7CRuqubI9vc8vqz3tZC/elf+JGv2CTfpLZX/CY/F6QNhUg16u4J
68Tu1Q/BX1o/4Ty1fq5EWcwZVZGpmRTWpFwWOJhT1Koss7Mt1rxpuxu+Gg4REeB+QaniqreIOoNG
uNWGJaRokDQXkJI0W3h0XpC5wEW1pcf9npoKbEP+ITkduhkkQJA07Jb/dgBigNyAoylz+EDEkNm7
LkEjVQDtPaTSLKhSN8u47JT8fQBmGVdIIgiJk0NMzBvKqSPLG6X2h8ucUmhOMW6BEVxMueOL8dpU
xB3Lv/ARzYshI2C3HKPjogmuhfCVz/17kIQx7VqsZLRvKoWu+t6mPO5K/YRfyfqouGxKjJ7uz7Aa
QCUIybFvGOPyJkjvq5lguLApSVjIjHq4sLxWjCIgfvUcSHGRRW96XgROPh4EYBRN8YzXLCy6cRWC
xWHZ07RTLkh2kW45e98hMwiJNDICqztutb3CRociETuoQWQWfUABIR/J/e9mXaMbnTCmUUkbKXoR
1HSVHJyDJqx6W7NJnWkzD0avmtohn2vyHb1X5K9WCfoxvg4Cf7kYpklJzMV8KwL64FY7plASyFJj
Cf8c1MNQNmTWSMVFXga2eDXqbcSsTfA/KGNllZj7CurESeg0S0CaYPr+WUWawawUCFqQAuw8eqf+
KlbU1Pj/164c27pfTz2QADlyePVD4NIf+N650BtZ6oWaH1CCvm5e0GHIQUmT/wNyfAf8kDbYFOf+
m704dVVe695159Ohb0Q1SXyjwaC8RWE1RLenQcL1hUyJ7fel3ygQhiI1k3qSv61Z7jQGMDp1rGus
GXD7j/2jF66qEy1Varxk00nydfi/ew4pKSULVjIk4alIv91CFj46LRSIDP1ZpUazg1nWFVr5oc4e
QybPA1XeE8HIchXXMXfyOqQ++TgNoweYGg1Z/WhA8r5w192bD8CW5Ac1am+sFK4+jzvqBqbS3gek
nFGTM/BK/aUxxVnH0Maks95keI4cT2uU7+nHy9vHx5ruYvvZSK+4YqhCn/++4yP92QGbTlmmLHRI
j0fp0S60EzD16udvvFun3zSZcMdOWsy8YsYPBEJKgBdUy0bkm8iTi2RQDlI/oyPIm2OVkFm/Zri7
3DJza09D3HGARQwRQGXjnlt6XBnbtGQgCaHgDOMEPkCPMe403e3sTo6k81ymsLdwNi57gCVwqZtn
lUFsUE0lKPdFY8Zbx4cN78LP4Q1Kg+vqx1RdV4NycD3o88OPU5t8OsugFUitxtEn2k6rMxJ0lHGM
Yy0T/icpjZzetCDxYwm/xK6Q3zdLE3pSpK8XAEzzugIL7+IuPrytZdfLGQT9c+zScA+IajFxEREX
keC+7TXsDSfjYAEX8buT+DO0duwgXT1Muy2m5VllEqBvvaKS/ikLUx7sX8MrS1AhEVeAPR0pDrA0
0fgopvQbUQJst+qntYW/eV3qA9JySIlxHpWocAUPBgCeFdG3Zgrv+Lm93CeAesQyKW2FrlM0B/NO
jYbKB3/wb6CFGNIyMhDFIF2KM0nSXaJFgPYDQ5FpDSV0+/0Q5cFp5ptU/H/zm2ymzE1lCn2m8KFj
G1RrIhNye0NH0rrVQg7CWsvjIt6oMcSwb5PiMGFBd5R6Kv1Sj8l62pdhfATsihzfoDWir+6JSver
tCCqqWiAHMUW0R2+FX/Ygena4tVcRIqoNHaZnS6g28m/Eqn8Wl59Hfx3xQw8wuKZMeUiNME/0taq
0zPdHfAws61CPsdH62l6QyiOtDk4Jhh0m3pWR/hMVuJQZaFNNzYc3VIGXDSyb8st+76J7b8Mc3ZO
pNF0DxbL/E76UG7TQVH6FUlu7anBVzRHjvOdtDzkoLLHNKiuh4iy/dLUEJ8mHEwBp/BPc0gxPeto
kuWtKVRCIB+XoR4W3M1VORaumuusIrqersRa5+3wzzjCtCOS2LPVG1IDMlxVeEqUEQVGgrB78cie
Oe8F/tLUfhhF8sASVEWdxvIWlBxPeZIYuiYuZnKQcj/oorZi60bwVjuBj5tthHVWSwCAjRantGOo
D7qzOA8CK1/lMsESnqZpnBSBnkglprgB04eNwSadJ9KHnQgkzMr6SJmXAEO33ytq/ORz+9og4TVh
UYqG5Vphu57ynCOKkv8+LzztGfwlisSwThlumIUsInr/5ZDGiU8CNIga199e1lFAjppadtYQbaKS
ZAyNYsfa74Yw/Q1nldh9at0b6wHX/t70XZVw3CX4XNtrXB4wHG85CKfFMNiIikOlCyi2RslFCoN3
Z1a3nmKkf9b4r1LszGlFEmbb1PhXdWiuS2kP6OQ+2BDF5Zboaa/4rQxTRvRxvuepG/5Q3+D1Ldz4
YIEVFkgPzx6leiiwfQ7qi85O3bywZ/54hHHBn2hn/E8QztG6NTWi3UcbqVM2Ql33UlQ2ss4I1osS
JTcKCKsOaeSe8jLiyAiDh2Gq7YIZmVhz5Uze4ip0z4wkTLbxKmImWwmrog66zpxhX+yT6CUBT9C5
jnQmqOx+1RQnisrlgHWyE4ctTKFXWrEIbNOPBb5l2eItlD02IuhjdZOAvKZn966MKMw/5RXQMuCP
MgP8re12w9cFOEzqXwMJt59w/FI3lQIo1CQj9YUXmKrpMWeUnA9QCXTcRfYQ3AtQAmsdL2ogvRHY
TsZTk+5Ysf9WOlJLXRpwP1RoC8hE78SwdqneldDf5q//Sn9u25Fmse4Ih7M3SgdxC6MJ4OEf0gIX
bjCTl2cI4/Sa8kLyqyWpYJRx9bV2uVxxs8PSy7nuUqoWfztQu2qGf0VjDFfpXfMVPYc/YO9E7qjC
lAuS2AgCpxoajLPUMuYx6jI5XrtYVF1BhfxcAbqayJEXLNGwA2ImNwwlUfmobBV++wsvhT0beFoK
BNakX+qB4G8E1hsQKs1QRugwaoiFS3oG28jmIvI1Cg9QCbS5th4K+Z6fqSNTGjSOnZt9XZbf0NbT
XBCysIq7ciPDfxDwW6ZYyT0GcnS6beCp3R6+18sRD4aR3EFAAaE2+DohuB0d7vIoZKxhIARDdIGO
EB9ejYwm8MrIv/6+sB/pPFVQaQ0rm9H2mkrlqAv+GK/IG5PS70NnDA3WCo6/xouDA3zKhl2f+b9S
/Nas/6LSh8dUZ+iVGa0AmppmqTmgdKmtqfwLQbNEyJA9Rh/5urcDTQh5bJSP0wnjXUElu7Up2xDL
xoHI1ltSHKngA90QfDn5a+KPpg+VBqUrAjJH6maLS0mo+rxObl8yJJ5KMckZaVIofTcvVZ0UMhoh
bRQTnkhKKsXIzmSzDBTfHzhjxIrqWLDuiJWbxBFCr4ED2gMS4Mx85plnY97lSyMOV0UOAPVwyIMj
GRz8TB0bH1vJKBplfk8qQ4pU55HS8RXc8JfPU3Kh850N5L+uqwLlDmuEeqOcEWCfst++66xBshN2
4zMUEDmv6GWkfNpkusw7VDghmp3KOxMTRsexvcXwA/oZScb7k29ouc5xeOkSsOHDgGNqH8S7C+3e
iVQSZOE6b3cxruuGHYUelMt2CsM72tvuWoBakNZQcZqYBpMqQLLh8wQ1Hk5YnVNHLdr4pILU7eoh
mIcfciXf4GwlZb4Q6yevUL8zAO66xk3bsjHOL646p3q/HAbOH8kO+ImUUMkW/yPTlNvlt3G3zpAr
yULtFhJdxzoOKaffPv9VNNMloDi8ChvcdhtXYkqY60DQwFG5BRh85CEWpyfBKc/glEYbP78sfNGL
w92URuxZZj0xz4knGLwkxdKrwSeTVodH5WmFWazUZUKlU42NxrbgMREjTEZpJFZJgHeOyGYwJ+8a
fAYetCG+En33tkjgjlTSlttZdygVyhThBkIszF4MZYamp12OPZnq/X7KwoHoGNwbIXUv4yFvzgRH
WylzUpdg8fXIQ0NfR2PRpobQ+9PkZwSpfa4iwXWQ5HfjLK0Bqs5+i2FpmiHWunMhcJc1CUvAa3Sn
BoRLeH7Jsf2vYmhNG9qPVhYI0+IgbUMsMmnsTK9J+S9zHXKN5HecAv14yA8tyGrLd+7+OipZ4p4M
IjCy0o1odGVNl+cQc2qiwAbsPXljtEeLwvzeeGCk/fKK1bFHrP2it1eL+Ci5kfyRqkW5P0KGH5YU
VpczUEJ/xCTmLBOF+k+pKu46YN4aUlolq1fqNo/gVKITYYQfC6n1t6QKImI5lh2/5xDiiV2FmaFq
rBu7g3n6EuwqOtpMMJ2QhmvynP2/4bmeqFR0IR7VSQ/ymymozfJU31wjj2fF6N99q5+D0rv4E0R0
wiN1iJPoBX+YY0hWlLbjgxhdapFydL6sdH5/eNEOeSlON8ep59sEysLoFEnOD7bCd5NQlnkjGZvq
k2hrWOX6lj+zrCcOYIp9WHoUDBDvgqGgodYPd0LBmZVDh6NrNyW6DUBqap1I6EeM9/x/CyclUwWz
GzCfgxdmuWVGAcNvo8fq6EKJnwiBpuNCY9If+I0zlYpAuHFlWUqSBYnK8X4JkLJrGLr9MTb8vpAj
ZFY026Sf6WTjmnNQL/9xdJlmfi+WjJU1uq8tq4ZhfoRxk73Pjz1eaCU39zjnFNUet3/5Q70Zn5Y2
MmxafPzDw0TEu/TnzvwS19A0vrD7E5rVT6ErVAXjnxICRWXlrH0khDepP1JSE/DGpk1A+1BPgfoO
Hu6S2zhFilb9CYkm0ui0ritcTINVNbSCUlhQXZ/Crn0TrdkDFgbIpvKO9uzPcftEf18txNqYw5yx
RPSu7iXO0R3NDjZM+X0+6kaPfoW2LD0DgaFFn4qcTr7aJ2VedMCUhRlv3sTi1/IqIRCGUPLmdmtB
+ugYGCoPrDWz4YjPk+x8vF9hKxvrfqWEoiZYJNFrVeX0313ryYi8X90XxHbbblw/Z+4HrM3drQl7
aaVl/a3DOpxrzXD/yhnahimNeZcSsEOhG9lhCUA5igdFFMDnLjGezDWX5mu9LhgO5JXzDD7o+HAD
We2z1AqsYN0K6VKYAK731DdW2qflQJG4gmoocGnRM8Xbbkh1IGZ+U/ntGuY94oYmOECURqbDntQx
/2c558md79VZ2yz98aArIgrMl2Ls6EZO0coeaNFapdBNhi0427al/jdYj3mph1PBOaQBtT9OYv2T
GTG4UMFtmHdCVmvrpF+d8LHv+iNmatB+hqtjdD2eEuT/OI0giFgcjysrfo57j1bAy+n+Z6Y9BlyA
w396x5+FE/6maPDo7M7QnChij3VDIgVvF4VUde+9j7kBHnoq5iZKFei5ekORMzuYrW2vsy2yVkXh
A538sBAlrt5sfZmkNdX763C1GyrJOVQ0171tmER+2smkXuV5EnSRnBIlWF9LqhGJD6TJhHd7lSyI
bkHxNGM7HHin+jmgCVI49YKVv3wF6WIenFMIvUJZbqrIPL/mpPg9iU0xOxlU6+mb/AE/8157CStY
iMBaG3FLv2Lxq0Otqo1jaLlpgHb6rLlcEmvncp9I7cxl+bdhixGdZ+N6lsDym4qWuLvKDs9NRDhJ
p33WptiHELwPg3elAKt5hY33i4ZYm7dcSPQPxTGfB6DY6f69B1g16hfFWcgJKMUA9iJNsfVfwliS
2n1LpDr5Fl9iHYejS8kzIxtYgInZQ/VOpQ2GiE/JvqhtyHIcnHsJ3uNkEZJzGkQBPctOz851z9rz
VUcUMSibQH35k1to1McyEvav2x4vrBZXKcjXqk/P+YcElWH4qW7cGt5yAejvVkgusAMImZCLRKOU
dH14i8/6xe2ylFN2XZC9d0N6VGMPNP/EqAx/RjwW6s5h59pYm6smRuUMQi5w+PqNLOWGMIpxCgk+
YiuwOWGSgZ141tIzPsrWT1vFCWI7Q64wtrIcX4nlIB1rk18iFHls51cJ3QUkGVBXQnrSL0FGZ5lh
uzU95khHnbz1DC8+lCLZ3zzodwNRdHFZVPtGLLpWA20aBPaMal2ni8ITn9EvGw4T9UapvEPP2S88
BWSSXk1aAzAIEs/lcATkCP4AIKSmpHUmukqBSD3h/o/UEzzzgpqgpkF7TzYKK/T5Vya00HhgTeKN
tCbs3u1IlYNKLgsUj5rWy8Iej4o/6Yp+IV9ZTp2Lqo4sH9Cd6rb4DVeLqADAeK0Kh17tUd8FitDT
MIcz2T6gfoetnp5TE8J0FTlZPofsiHjRH6GZg3w9rC+vLRZNonkevakrcJ9r6AIR4phWu7IyzC/Z
S7q2Y9sw9tb6t3TWqPaFGFxDffKvuEsryEL9+z8DfTL6EqgyghRHogzxW6ee/BNqeXvEDB3LPlx3
vyYRYiPsgYGXFttnjmQJc825Mfyi7E0K828d2Cma21AOYgw20c4W5RtsfAGUPa5UbczdvYhpOAZx
RlFR84hhJibTy88DpKVSXT4h6gaQQ9XuK1qnlsjbchVnc1cELq8o2+la4sX60DXwuj5JBhw2Cvv0
n92yCdg9A2Oevl80JsIZa6Ghe3+jwhayP25sEtN452olDRgtsE3FvgiJx2buCfgTL59KII9MbiPl
TQuVF8+4VVqk9eB3jk/nJ+T+mrSwIJ+nc07NL7lN39Ap5APlDLanuyHbxi9Lqe2iiwD4fEqIoEe7
9+ACx9VAox6Q3SU45K74o5v0pM2+NcHS1ZAjxR3R8eM0ONJ0hjRXU7pCyQY0Cv1R19tHbea1sAxM
493NPRjzTHIbd3w1V2wnVcyBib4yrKKQVt6GXAPD19caY55e2sV4ONwnB7kVdusGuM2fZwSVVMoe
jfl06DRRN/4QxkzJFhY3zjdMokmSdOZEgcFLSfmr25qkZaad4+90Qq6dX0DX1strqjjRB15mYnuW
WRCdDbb96zkYL6NtAymqwrWAGDyPrwuj8Xh4j6RExDQwq0VlZvL7F4GzAPJDFt+tIg3rSD15VaoY
aesV/87dt0OSFb/lTUMe1ntum7nkyap9+aK+uiyv3LmlNzQGW+jFso81tK/YlYz9mnSVQ+Liw6xg
4ZZcRBbwrtGZIU5SjQmSCP7RtSthcr2bizznr8r/jfZQKs0/Yhp7reZrrEU7i6haNNVI/xXSNyQb
Runj283jIGF+Cye1Ct02HjlqTqk5nbEpTpM+zYOpdV//eYOKCDNYgPfee6i5+uemOmz6gUmbf0Ka
Erni8D/c+zULPH9uhqGfR2Yf/xZDh1tNruznJ96IXrvwS2caGPn9CJbZ0eY9wqBuRtTG56jPoL75
GPLeU1blyootzcxyWuW/cF9Rm/pkyYDqS1YT4jgXx2OqceHeDr4A79yt3FIald2RDrANiB64J4h3
jRzNBSU+Ni+tLMiq0EQaIs3zkeeydNItEhr7hy9PY0zWAYETisVFeQM4CYscs6VslnMUsqEi7njg
6QiNomqRVkGntRDvQ7ZCsAA2znk/T2XGLdPk+TafmsnGSn6n/QfKQWmrbzDpVTzlvNvOqXpvMutb
hS3HAZFi+5IsmYnGhqoXR8socZt6T7r3OtOwbZHKpKdzQJW1mxGN/FSTlJgCS6+GqXdpxXen1SOr
YHRVnuzvP5fz+NT5kuC+OkGF5SvJty6Cn3Ubzh1Ti0J7MhPaMOXX6tzBzcFRn4zx2Iel2lcKtz5U
7BtmIQh9M0Myw8ncIj5miAbQuYK2L9jTD6XFvkL3I6Q050wwqW7fYnLwWoGJ6ZaUI3Z028XcR+GB
E2kmsHW/WoyNHKTxqXHjklHZ26OT+12ChO/IDSGAgBRdH7RtC8MkGGOTjP1ktDQLFqtmz7/R8Mup
ZckpO9eBsgbQs8imLOGuA4uYlhA3Nb/wlqiwIcOL7CKvOk/arUgVNmzdndIpyVJDe+ivF+4SthaD
5q62mahuF753yLcsUafIU2giEUWgLiUtoShJjIjpunBuOIWRpKDmc3CCOQ3lzzIS24P99PZ/IW7U
hzKIQRQh0cqFeSaaQGq2h8mMm4rtXg9g2IXl1mdfq39lyNlniYF5G+0IQoLVp9inh4uSuhW7pk8l
9uTOlahgddifzvPtx6ra3O6BOvMesPnNP4QsZWcaSmp3Lbsj9ne9ulJ/I9fa2iTd4y14dGi2NysU
WivaK4mZEC3e+8vjOtScFXOIzjUIsVGfwfa6CRDTx7gd5NsNEQupbpl2bYqG4gYchVifU2F3THVM
c6BCrvvK7Q9PeQS6Tdv4C87wL+ihnSOmv5gq2FxERzaTIrlPZOGtUnogOQo5R6RLuyXhxI9zT4d4
Cxm6vB2IGm5jb5+XBPkQlA4TQMedPJsV0rUdeoo/6m6ivZfZW1rW1PgUVFVH9fQXnzBO7+MVE9Ad
/bOMBLdqQt4dahuW13YcWYuPsFrnqKZW744o/8HdSEOcfsnobflo4dMygJFP5xXpkAcWV8aFehVW
i/8lxSV3/faOhteQdjZmZX5XP6V8oSHqgtaLYrGPYA8GlWOoH4LYxW08JAjuOE/Kz/yBnMr7Y6K/
+EPhDoYqEw3zSYQjG/1rwCCKZsLMJkeZBAd4522LaQMEOWfwDTv7C06khftLnA4NpYDk9j4z1W2t
ZK2YnreHdkQxHbPqBR6wVmecG0l0Ps/O++M88kzY8NXTn/vUVeWwN9ebqyjVwEiwLnJN2zS854k4
uHeAJ78QD8mTJOHOaRmkMGR3yS+Y02aB4aww0abBia4ykJ6RWHWQQCp7a+NQSQ05XlJ6a7zb2cHn
kz5A9zrS+MrPut63YXRUJphrrKj98+jGI0qWrJvemxjWv7ZWJSeMz/OWKRv5wSgNuiBwW3Pgb1p3
qVa6bZpYfZLm85meHf0NIMR/2oo2oM7i8+o3Hfmbvk3bDiUNkwmSjT13UUSM4ZB/B8HzCiPMcHu5
5lvr+GxmsV/mtmq5jhKCIBpDoY1+/9eEWvjAAK+12KuBkhwoMwOi4E0NvbMLcWqxytj+vIZhydEK
oXFPfnXtKfsUdzzI0PeiarAMp0Ad1AE0Lx8V55puISEDpUmFe9akEw9vslLwtfl35vrRAAp8FcBr
ZJy2BtReYNB5zVy2TKdSAH1llv3fATonSwZzXQnfFKbMJz0OXbtLJ3ZzvKWDFV5SXo1IYNSC0tEx
Fzw1DVbIO8oIBs55rZKdI/nHyNIF1JD0iDdIhpMT4l9JURGHGSYxceLPzFc8zQLYphjRzK75nIyO
GeYCnk4rf5IY1fkNNGLbfX7DRekkQsqyp/sn8SLefEOtQ1IeBdX4G6+vS+XQJ6FoXoJfDl7Cfs2r
Y1t+Zyx6eiTGZbC17GP0x2kBh7P9Q7iq0OytjBrj7FSgdJxG7lRs3STtClMKufprAGoeb2g6B9Le
hkyMLr+9/gvBB82G10aQreS2TU3iMzsXRD4qheZE2luyUnWJkBjONIXjFBtgVtnwKXJUY9ViNGpy
Qay7XQkxAvNBRep2LgzL9WEZ71YLhKZq1QXcFussitKhvU3HwHvnQ5VTdTeWmp3Zi9TfRcFvrGmf
g8X6XT3tAbX2KOlOEcLKd9GspPvmLVzWP9O9nSAvbvxe1BheGbJpS2jUd0msn7ZitAWSRHjVz4sC
8vSyYrPl9oVeetOUp60rhcfODXJZTp+BkSJfSvv3O/RJ4ZvLOgUynWYDdFRnX+79SMRn9bFYb+Lh
VdWgAvPO3jk+FAyYIy2//Rxj19QFPegkPKRxxrlvl4hmC4pbuSubU71TVY5fpBvVPYWYgpzSpFPD
uiULpDpYgLAYv5NfURPalAPJDUcf6k9J5pbwmNi8v3Ohz0sjgbXInApiy5IlhL/dxmGXgH1Rk5E8
YW2ifpXAQCdfDoBoYH1o3uPuvHz+80KlwvL+XeQhmGGcbdiTXqDDBtbKRGYU0UvR9OAfmUA4MzSS
aBY5s7ef0AedDr7c6R4HZJEG+YLzF+ZTruErwnLjofk4AfkxeoPuvuudETjldPOqnlen27q9Ybp5
FqvAC0WiGVLvJS2RTmH8IGhyqT+0gMXenEEXukpAoZuwDyi0p2rNO3/KmUpma2L/hwwLu3WepiL0
BfqFqWfjMMN/rqP+DQdAMjQMU84iNgdQqpXEhHKmrGoQxjFvM1eiqVKZlW84l1IOlpBYSHbey/W0
k2ZZ0fnRW7DO3Rl6obJNiG0HVd3+wpZkjdxVZ6nBA1YLiEdPC1CYqbzbR0bruE43fZ0viX4huncE
4ehhkYfKzNPxoP4jlAe8j+PY7rQqSpbxXrC58dWLkR/MiCwTAdXfFuSTGEhNrpTIdCdmIit6pwzk
DIqQMrARGIwbnhUdhKscE/RUrgccH9DbJGupSiYx7yF1kba4twRo3mqlV31QdanVLv3lV+gs1qru
68rb1eQUnwdYTMzNW0KD83+UpNlHY00nSge4iTzPAzTWxA6DL3zpsz06O1XQOjxcR48SgFBEQTyl
hLTY49gRG2+Sn8bZZrrGRwiVX+nci7vPhO8Nwojjx9oKVypr/Czg8Gk/wD0hj6XFkCwzqCtKjsBK
OvO6xUtmhddSSfSmt7xegOP5MpjEY+7rPsGTi+Unw0/VWMinryP3sYqjGL0OUBb3hXcqy84oqBPz
p6S7JRDmXToZf+seWored3KpwoNsxd9+Anm0X+l6EbUTXl+qCKNzp+crG5N2+UQWJ52vmxZcN185
LGgVLB9MehQZ5OA0XhNSSAwavtftB0KVpteBrUTL11kZ6+5CsQwEPVJlkkdFg0gXy5xYYLG5ParL
FjN+pxbJ9UXnGPkhPxALtgAWqQ5BFv+NCRS0WC4CftjxA/ighiRW8lreCRh5fP71ICc1EV3nb26g
s//tENJOfnTyxfQQEC/oAQxQFHEVWjojwhUoxT84omwYQjBJ+Rcos5P3h8poiSgGfLBNiFclIg0p
i1jYyd8qZAtirO4btOv3+tuirOJzReWfZ0hhMwlUv102lc3lITL6bO8VNlJuLxbHErPBhrK5bCXa
n/J0LupRNNm57zfY3H/jqx61MRdMmQuJYDiqQ+9H9CDaa4GnzUooOyTIcWFgXS6a0CXVhw9ELbQW
uBG5JzTZPyIB07L66KKNCAusZGdkxyvkgoCSRDpn2oXXtFC905qca4eydoF9vWZKiY5Xf/xIF2Bh
8TJlERr9ERCbvDwvR7qm4ZiOS5jyHcr5hiZjW9rLKFcUHuy8VvcrZAKdol+T4I/ePKBwthSjbHsy
fvOo+PlIIfnSyOHhWQBhkZnWQ3a5UOrlaft5UEPw+pui9Dit0CAbY5fQoBiroTI8aXvGTqAJQa/V
h68utaVb6Ck4m0bDX4GYU56O87bua9SLqusomna7zXEISmNf9rv5NcsFR15GHODWSxwzh6vSGqch
WzRrnFLaszPq5afR8c2DTtxpTc8LaUo0xrB93aoyE3MOvSzSK4Z7IWCDLSBDyXOL702d6GyKvvVZ
n9Lh5u5xJU5lmP347+AElm8bZl97vSv34hcPDuvaTKwyF6Mm2TFueI+NfX+Qibmj1RfmCmnt54hJ
4yX8vUSQTdJgv5JgjfQB5RVA9jfMSfrYKgOIczFCKeTi4W0Zc2pfnW16jYrVePj9Rydt7u0JiAxG
LeYjWIavKO67nTCN6VRi2hAqKZvYhBwHSXCTp2SjPTZyeFpiSRW8DDEMLb3hpPLrx4UhJOlvHm91
0iVgzQSmRlSDxSo2lZCRDAZ1n1PaIQTIJEhzsjaa46koAWTZ37m4Y0JLGtIuECHsWiCrpKzccMnI
NBptgRyIACr1DuCcmEboANSKchkx4QUo4h0EGuth8qFpqY7c7jpBBU/FU3KDVwLQEBFsXEc8GTyb
lF0RKnWv9VtlrpxiSEWespfzXWf0RgCroKtQUh2s/hF3PkTKewiwhqFYbu/XB95gGRPlhQhcOBh2
QU+yjYCLXYVnOPCoHPQbtAZGolvTlL/GKiHkNN5VllyFyUFb8raRemtsf41V9VuzTerqu1l4txmj
OgIYGOeWSmIIw/k2TQxE1+qLeXr9K+Pc+vEFP0pjVjN2a/ujDKmVdjSyf0mEjNzfzFmXLENKuhsE
8t3eFyFtWxMWBehI6LWK+EAZxyijghUTBjyMYaP/jCYt2SHZ37FtOjIGmEQ9t9Abf1Y26KB6M+bu
El+mmFoNphC1tDhqy8QxQ1nrmdx0wwequ5DhBzi4P5ddELJ5aTz/YaLH0mORcuY1F3TdO8PUq5D2
I/vUZDXDNyAbDttSTo/po52QJPOk3oHjobJxe0Oeq2OGIhrVjVseWQkKfqjwW1aVyRO/7GWvEPS5
3BKrG5vmPepvZRWpNs25EpUCmhPa4bFWSXLIY8d6PVR+mY5bCjRY9efGRH2rPJmpYfen8Oq78vf9
mnR6+Wmif+3zVM9QGXHscwImwyzaCauG7+W95dHa7H6NmTvfyWqGf5jIRO0ulOIfGfzMXbsIYvpt
D593PXbtJQrrmx3EMrL2czsLHFWrkqG/Gz54qkQcGhsE8nLr7IuE4VbFUxRGUy3smyIg7L4qXFgJ
Eh4v9Kv3q4sxE1vCVUhxHkG/p+2eFDw7Q4Q9SLu6QVfkMUNn4zfS1rknyLBL7BTih2ldtL8bx8R3
BBwvyEM8CoJL2ulKNlKA/bqF7KB4qfQoNf7J6ttf64auooMVGveUCMIOm2JHsIV+sNkuDvYghlFx
bFMJfDJraYv3/nITQY0zUXRy71mkjT+RK7BJIO13bQzePxnPDT7rf1pKzm4xtQGtGx/xmhXuJN80
ErCnq4X5TlHYhl3Mxgg4Den0X9oyJXRWfmWo0U5zthgFDu0/Bt87uB7rKnEkXfDFuCrBMTd4fhUT
64LjH9jSKBtwHblJKsyzkTAh34N/m6NA2MuRZFtnEedBPEO/R3kxIF9fQcxWe0SrTY88QJVEyYds
k4ktZnkpddazuu/h+ps5/sFlza6rPT+JurJe2L+NFyLrA+dSscguHVb829y0fOSqTdaUxK3sKQQo
R+f9VkxI0vK3C/rn2wti0nYfCeUTL+g9b8SPkLZNcnUk69IzzRkqpGIZhyln3v+un2t9Fn46kanz
qeTdKutA2gyPGYOMtUqPpNWvjdsB2jAitXT6uxidC9tUEfxVwLhSTYUdJPgpyXE0UvcT44oFgodf
qIWwvN7do3ZjRYeyLZCY2jODpCeoJcDm4zBx9ZBAfPeNFG/ZxXXh4qscrpE0yhZNdoF8nUixKfHa
rMUoG0UbvZzqygpZyx4y1D1AeTtdzA5nt7k9YAK8u1zPDertQbrgycF+oldKqabbOSSpwuRbXmDu
0KoEuOP00pLB579Au8FJvh/OLHjSGRooLlnAzJMdbVTPr3CPGOyf5+1gGpgxizRGILPwea9sV3bj
rs5EZeKIebuCh1EBGSvKpHwPBAX0/cTzxsnwrertzFlLSk15XPr/6Iv2nCg1A8+eP8anAi3ZO1r/
GASTGibeesgkkVfqWOO+pPftd+Bsw0iE2xDVXA4HwITRjsKT62Vp1o/son/Nhgajih3EITa07L62
eN7S3CAiqjPtMxc1WFfGjTpPJiR38fPm00Dm7fXm5OJjX2YapRaJuKgBmEtkSYZb/TSfDLHGoyEX
AQ1YFMAD9CSo5wQ0YR7fg+AJTAsfqVbflgB+BsAmVU5nnvKB3IHYeraIm5BKUlyhG3IW4M9OgJ6K
qQybyivmL0gEBD8RqCcSrI82JmMgWfUWTKYlzu6ggPv4bIavmecgX+B6cWf1BaC6mSH9sRVhOg+K
Y+ehG+tVFqBDXyZkP7zybAjgS/H/uTnvbyAC3UOkt3X166hVaFyHdl+hlOYNZt4oWi0rsjTx4jJ2
RreBWyR5pbKQ/OMkA77Dp/F3wCrmxs4+GPVVym6kXhyh4xQ7zzY7bO2SjU7l1IqvdJ/1nxlrd14c
TGW8SGknO2/i/7b/xcOhn1zZ83KeaJemijJi7+HhZG8KEavKOSoAdfgx5GVJHBBdrVr07BSis+u/
dWEFF1NokXlW35EKqZdLAOXHEjFgCDd0NrW9qmABWIdIHFVbg+Zz3mMIdcJarJVANmTHf73BIiEq
GOy1FM+GTs+wOgjd4U3BjhMRTN8+hYHX7ky72l6JIGbSoP4p/Kyxg9eSkwcVrk41DVuwKbdZoj1v
Z1mewXbKPvHkOOeqHkQS4eNxRcTlDdAZaGEpPZLl0kksXQeQEghqKdojxgCg9SWCHhIGH0ScV3Xw
GF2xHM83nYeHzWjMK0nzX/DUnJfYIt87ze1xByssi8MUT8+0pKxWHR9SS3iKFODtMLsiBFRGhhJS
z7OrtySn71bIZC/+wYalW/pHl60LTZKMwmsgM0OIruLQOYlErilg6fiTT7yy4iHE2r33WCEzIltd
Hi6nJezRlvSKuUGKMTVUwLx5IIpDhaE82MP/lSelBQIlKubmE2ureyPMuDPHXSNUHjtqyPW1RNek
zdD25XFBflBs/5qfYmPK1JaYVpd5GMKn5JuYrlHJ5Jdx9BpLEaBeXPUYMAafI2r0+iDGtX+Ycl7E
CKd43XnHtEhq4hoaZo8SfvhNk+l5Hd8ZQPGA8vcnNPKitAR+8TsTf2V9YNaPGugcFkP1GjMa1ddd
wBjgey9SxlbdbVyrhzomXl6rfdWMFaOur9zTnDKa0JDNZ3rPlU3YLTedfzqSl1fWdWaiu+EpKvFR
XPaS+PyOFkkKePZPYq9Pm4eIxxq1GBukdr6aXV34dHmnOFs44oWnkbIrJiXQtaIAWG1PKP8qAlY7
5O5wRc3lqmrHGVGuhKIfK0Rmtvh0JyKf4WV/ZLnFnnVHXboDCnbq6+aMjTwUiWIWpfDwm77+C973
eFER2RJaqcm+nXthQWMcmWamIJaMhfnQgNcj24EWhapKRSq43eT3ZOAAZ75BglwwwCmfo5OW07sB
r+rQds/MpWtzhX3cWt7FIzV6PYKv6huRlPg1j/lZtB7muwma7+Tede2jpBpFSkG9Sbsn8qErHCLU
5xQ/a6I+U9V9O2eXogzA/77vWnn1hDWU8AR6YaEw8ZCGtr9iNxYpGoiiIsi2f3qvva8nZCdDpHur
iZIOYJb87OuU5P/c3oXJfQZ1cKxYNOIUlwKfujggFumNQKjUzxhrv2eraq+o/u8lBrOb8SPuH1bk
bdsSXpvAnsUpY7alWs5QiI+2aLiTGzuqrdp3lPQ3LLBR+MaIBsnbbPs+ZHjDTGyPRd2KZhyABGzE
JPFLu0ifgp7oWyJXbukuGRRVeIsiDJcGozdNzRGANe0BWQwW0U88gwWCNR1gwD1Y4aOhVEldq57C
7qkktr7KGsJdj2xI+Tj6/OyfEoIuDhveDFx8wbbHpK8kYWf84juJoJPW1tQloLeVJcszdWE66QQJ
h/VxhVcmHkIju1n/wvsW2hbogpgWAJ4RO+9mVi/yS7HyHFc/NDxD/pustbWHJ0L9MXF3dHJYAQG1
/V/0J2M0R0UAJGVNSFD6K20iiQv6xHULGtZye8AWoXfQNpd9jOmj2hoWNiLfhSJQVZQgkUo65peD
SCgdU+/XhBA/HpkOfcFpyY2Ll7jI/9JlQiFuyWm2Bwk4GFhdH9k08TnOlv5Cv2XfxfmxjToW2QEM
y1R4w6sqBDEHeAJiuQdlfKVozHD9+Vxuq+0oVONvR5Sq3NNAzImVW4v2cdu+wH+BipL86wO4Zh3x
KkvfwFfBIzCsndDRjJwFkR4mkZLvzKK/ogyvikNC2fvhI46PjgjU7aJVIaaOybLo9U5uuR+/acuE
KyjTzy8Ziza7qjEiqgLxKdk6D2Dl93Xs4FNycn9eiSKnKRUeGNfwVs89zI8EgYuwOxIhmKljprqG
dz2T4yNbJsf0zIb3TH8r4RnclTy15dAa+7lVZAzEXKuCbB8dVTLDfU13aRVN04CNSAzZcjsoEqiy
2kephqTRq4/JPPf75lrqtsum5/hlhKWnhDVaxkz/NNbzMg7fn21VQ82STDdZzxO27a1lO/2vKwEc
7KZcbRvumty8VY8eTZ/zKMaMruMsZCZfigBUXMHdC9E2ODj/3IZ/7E+Nzhf/U5j/ic5McM+8i2XY
p+TBq0Awu8nd/ISqSeDObMEXSGy79EAEd/DO5X2d2LmzmrjOfdh2hGfDc/vjZMcjrwSapCx/lVeq
Xp8GN0UMQIPj0PxpX6ZZbog5kIPn11aDuuDctp12Z3G/fJbKOFTFOYKAkrfB5bnoc3nERSfS80In
cHYRA7M6Q3vWX6cHs1RcX4fdSymL0zq2qhV5/qmXghRFQ31tNGAyw9zI9da5FRSBMJmw3fpqtb+1
ZvtZFOP4J71YCi0ZsqfPKnl0X07tdzKMgq7RBHfjIM4//LxmATP7DS4BfhLjMOfqBD1upzwAmdPO
Q61ZD62N1idzhFAma/WPYTuqa8ox5qa+XOM5vraupXCB8VZ1U5Xt5uk9hNsNyWVwe6dv/8rrzmfi
OWxKMbzEdavZQ0XS6QnSWs7Me+XjORqAHFdIjrqyrfUuj+cwO6FOKsFjXzVfTJTiB9TAij0SJenk
jcU52Hy7cQxPQnEPb+7pkeVe5QJziTiLoiv7LvTSegXZYDTvDU//JVeUYeYziSA40iSbsVsEbCCs
nYXnQQZVpOoFnNt4GD8mUSN+wOhsPZEZK9mriT+tZBFID9mQ0rk/GWsAyV6dWJFigRRcc+QAI2h0
5Kkh9Hfxynv5pwOfk9YOA7TWa8thzpT8NbAq2FDfijDYoPnol1r/cT9CNhhgDnXtPCYhtkFOlsqN
BdjUslT/Hcb+ll7MFseJv+sVh/YuGP+zxMDoAhfXpJ1oKpbpJehpxXxEdPbvEULffvf3TIdVTmSC
vbsAk3d9+QZlZReRXgFIVABfguL0xDpTrkSOsSlwKfujHSO0wPj08S7VFtmgWFluOS4i1/Qk3EHh
GZEzL5xCy3pulHs6wL2wbUAjUZS2uxoARUpp++XHL3u/HAba0/o8/pZVvGC2ARSHKXdhB0pIGSX1
wUH2ehx+oiwx1s7/Owe2pPH+iow/KrwnWDJEiaDODz9bI0OwBuvjHZXIFStNdmI1ZDbabZQJ8oTC
ZmR6/5SElGyIW4Ht4bMvA0jSdjxmaMCIsfyHtIqGM+wfaUwTxtiFI45OBATdTiDU2W7XZSUcPkYR
bLTLd8oyrrx2sp6PEg8pd+F80Wm5hAFXjcmPY7n6WsvVOvkq0saU7fjfvqYNzUeNL4TweIJvRJ4b
ECM37dA71clHqN3hTCkFB/q9qDAYmpVagsTQOeRPtb2QY+3BEW0EHcbiwEtfQzvUJx5PcKVDGHI5
WolHL31COTRtOLAAxRGYyfBJIUUewCI/gmqs6AnBxNiFJdEEBRFm5OLGgxmbqJA4yDlWytgJSQL+
nyIDtbHt6SBxRpj3h3UDzGc719h4ytGnyHHX2Z7Pvy2q4/Q/bhVNPU8zcA9px+8rJSetZAhQMKzh
bNmSKbSuCvuOwMmkdfpwvaDAjLaM8UHuvtNspB0Rn2FzVlUDPvvnVd2p4BnQZmJsOv6fKxNfpm+1
dqFhI7IC6BHoNhS4nUg+3dgMgpTz7RMyuXVbP1OXoTvT1pSqLNo7fvEnkFFbX+afgZ1PrmUSYtjg
z/g7o5XesdUjFhkKC69rSwrRNFfkKJI7w8CQezVqAOGT70EaNSas+riHFhFK4TGkcbf5QrbAhJQ3
WeQXMoTTSPpE/QJmM+h6vOOS+WCr0VTZajZfoRpDPeJHH3+dwculZy2ntxq3P7JsocIdVY/xfH/Z
AVmdTcURz2DeYiY0HzFgq6wF8qxzp8UY5MslGcNHmiAhP8P+vpTsgSU1ZDMZrOd6UTJj0123iPKR
1TLH58ABqLfWujaC2g8081S3pQNkRM91KbtPv4kZkNsQRUYcD/Eeyi/VH6Un2xRhd0nCvbbh4n25
7Jxf1jvjr6e8jUoD4qRQnwmOYdBhkEHnOUXrE8sArazm9llkBfP19pBnMi9ckOjPRNNuVRQKh45f
DTWUUN22WN8GQ0cBqBsqxnhHG6rbxT8hsRnCPhPQ+Ccl402zF4FT7VXdxVwqAb7JkybfrZSaNK8G
ucPDnNpqz2dENEjxaxLHlbyhXWf7EdRK1HjsvCh+eT7Fytt2jE/GkpgwMkubkO1ypo0w86VT/pgW
u+w4CWggg3vmq84pY4hYZMYR59csztOEjv9UfZxRXEx02IWbjIE+xLWYXUdbEJ8l3gI+3l3jwmvv
Ciyob+MxPqNz5ALvTm+n6HMrZz47dYwM26kY1djy3JmQnZ/5XFQkODC3A5MurHYg6Fibdc5nRtx8
JBOcyCAoliIGiamNfj7xH+V72mF0wG7AcSpk2+VHKGw8Dx52GQ+tBMFuejDkbsKB5y32V0cGQhFD
4TSx3Pi2J3XiEbLOiKI+nsNrruio/RtB5Pc5TJxk7uD/Jt7+PkQMh5YdEaGbGwOd/lWIvDRc0pMa
XG8uQ1YaRhmgYEpHZZBFAcCYsxNEYiiTd6klDyyFzCufRvyApFP8Vq47vvKRbCibdkGRusyMkuiS
KX0vgFnKYUV47q8uomKc/WNuOSqEAH6MLy8vhIUTwntWac4aI6BJm6eTG9J7zoEvVWv1u654qvmx
yfa/+InBaiqckrUZ3HBHI399S5akurPiZOFoscGkQsBEvtmYZJkUykiAWfbyqb9nydlTRF5CAnjq
l21QpmHMpCybVHC/e+bWysgrl9Y+kjb7FtO6rQPMpwc7Jo7VVBnyMyP5PfTW3BFkpstGrnYFOPLC
hvjx69rkFomr5b8bGCdkJFG8yjSLcKcOQiop8X5ewwWteIQsTtw3zvXIySy+oz82P22DSXuHXG5S
iEytXIwH05Mw5mHWwR2caif+R3tvexjqrccYhbdMVeX5yvhj6M4ZLCkSjPWdNhcDi0tEgTfZro6E
RILf5pGSLzB9mi/u1aMyZA8R3+PkJkQn+k/53vHV9tV4FIlLzXRU3fRS7TLhXxxKJaZz+T/wapZZ
IqH2WUKpfC2GfIu6Ekcu/PP8ANurytXYkqMt2Z3I8u8Fmi4tOc4iYR5pFqCAZWVQmW9Dz5ZWZnyr
4Jkvd3WpkTRdkc10uITte2mSmB/U21eidIf+S6W6I3EuSi/hbMeCyfu1vkOeTys3kTU1AhoJ1Rjq
gw9XHJlPjd2lkVYWkn+G3bFu9T+euy4fWDSqEWXfqcf28OFc6KzDcqHSjEyjKpZIj1ckx6lNET7F
wM/mocvJSvelXvttbo39T9ma/iirA5DFxQueRL9S3Q4dO2NaN7gTEXV0cv5ad44b+ZIOTvI9xFjE
xppmWOSMnGi9JsVewMio03uLwDqWNTlPEVCifLk5zfFcRakn5G1SfWiiUT0d7RjHuHrbk9Lu19C/
/ENitjXiNYijvWh1Qm10lxVoa0PiHvGAWMMulOhW6mUeqULiJ84mGi9P9NRyBUfvZUugA4oBYQRZ
C9uJKnFSwGoZ6OVpC+tFFTc1WxsjVzSgc/5SQQXzUHb70rthF0uHMxCHaA9XUgHPrWduQQxo2xPq
hVq8WZ0UMHHTa/k3IU/eZ4Y09fLMyzI28rA0r3IMX3F+nb2Z7QpxTcQfKlFicIoxtDiXcjC1aL+U
oqmuao2ZSHyjBOlozXZxmHZerweAmNfbc5rP2zHaJPndPV6QS9v8fOexNY2MzsnT2j7lpesCNWHJ
T1I5bMhuyJ2dLA+JwSeepGQ3LhLtSrp7pW/cpqd7ZXigwacNfdi28Bp98zaDeK+2WrYyAFVND3yz
HvxbQw5ey0dl7nJTnlXF2YdgJj2KGsW+kNhM8rzgQM+XMfmjZasheIp8ZJgZ0RQPxCbCSaaj+4jL
iUJcOdIh0tNk2aqUzP+UH2FB1jq0kC9W4ez+2y9UvxCCdGFPVh8DoAQ5faiqW7dsCbtGFN8huayj
1nPpkmRKNz7fNu79RRqifuT0AUsGc1GdX7LdJECGaGPRW/8hT3CuLcuh6yvE72yIpCaa2a1Q5eA9
e182/aOcgX6b3qOP9uhfPIvEO/Opq3fTOjwuW5QtCCSzyu94SouKgtePBYRd5OKl2yybvsYtnAGe
Y07v9q4SuNsNMVyc/M14vk3QGBALRgHKRy/kME3fEWpfYDMGhnWHs45BrvImEO4YZbgajHNZgaXx
wASBPGr7uRHZKI+fuGXS9k7iakzKH5a8+FkcnfUxkxBLJWZB3bWt0KqinaVQw7+97rowb4zOwRt/
MKDFJ+1NuZ+3P/IMjqMFNFt27ih8HrAs6jBRKtO9Hk5G/tzVMchpcO/2NIjd7WOdmFMy5r212ON/
rFv75xlA4nsF98uwtVwj0slFIC96Mu+wk3sNcjlZuLakFntaUPK2x1pZj4Ev29FQuj0e3IRLMT2l
pX2gE062gcMxW9NEI4W+dDnEPTYU6FiYteswR8I+9o4ybu+CIcjMH2sF3Lb0n+h+UFRJ9qK3PNl2
bVm1ckWXRYtxoTsi8AGVuX6yJC60JTQ2qG/PR7osx6swos2x84woJeACGz9VAHpHHFZ9WlfcQdwz
CHoFLbiyR8cMgF0N5ef1nzBihv36mU2fuWiJ2sb79dZb7YwJXgvLrzyGoibho6rnvXT0JDPIkDZB
k7OlsSMjcpZiJe/I+zrPjF3DbNExaoFYU5hrejOwXelw7K/zMKolPrxY7yoAkb/XtjF76NN9T1WV
7frJtDs5kMUsKKem/b1lQOWmfO+85+AAZT+Gof5zXzswzjWAuUJeQwaqBgw/vQzR2On2MOTjFGcR
sBbtcMy6KPmZRyTQe+nXP4E0ae5CXLJ0Timr3PyqoC/y+8O9wjR7y1N/53MTL5F8mrtC2Sc3vqdU
2s5O8BT3Jh8eMY+ZnBh+cR7pqjjU9vfBLv2N2zA6PlSAqf376LSzoSxVuWI0JW3fe5FWWKG0THCC
MiMGhpflnwbXFTPcrkciFYU3V35EM9XGPBtavBm6u9IprtLe6hUvmzOqvW9qYZi/Rl7/PP20SIIy
hZJDxGTgqKoKxkdSdC4Earr9cKc/3bCG1v23MBe+1UwaUTsIznTYK2ROGr22Ikm0/Ubq7IRAjZC/
PPlShGo0OOZc6CiMGa1heyfib2Ht84sj2XFSHNipgTl94pITcderfXquoscLL8Q1YzLWN6PPvCIv
rKU2zjrXY9hpP90gs8SDyVIIhtoSfnQ8CGb8+hgfV8vxSzLPFeVGdWH1ataJidKToHNsH+bSEX0A
HtQtXO5J8KIrvxm4t1K1wtq/0jhHiWhGx99qoQpXKS/b6w7xdWYmVdt7c0ZPJU4KnrLbHSHA+iMD
WGJD2nhHaj2WkFRz59fhnkJBYOTaTpJ1VBc5K461Xi2PxAYp0UTz6rvnR5Lupu8gEhQxq6HhtdzE
4qo8R01CRUWqLmf0b2vyCI8ilnAMgI5HcbLIC4sUNDQBQIa/H9BFbqNVPvVncs2yK07tmuddPq59
UzNi93bwFuT7iAkYKzN7whGmrastn0iObExWQCLSTxEoIW9rLlcdHIGqOP9ksLo9gp6Xu6sNKeIV
LDHdeW7vLSidFBHryb2UojHwXxIl5xBYrUK3lgqYTfthGftdlATgxZHRgs5lFId1DHTsU2QTJ6zs
T7Jav725lziPbK5CE7Pz/nNtkyJ9LbMZfIg/vrGBREfocYVjRWK0BLbPKa2K4xlAccNgWLE6ofJ1
wADEvLEN93qiMYZ1r4Kjv1QwQai4HcwnEhGRAaSVBxWmvbFpxMzWyoqebU9cGuxhsHINAnOxdn2t
gCYYZOibf54eRCB9KtThCD2F0LuLwhd2yxs7NxM+QCQktnPJxubmE/Ci8UzAH7bMZCsEzokvN2D6
XIVwrwXeFH1cWc/2Dcn5Cf58e93yI0hOZPt8rQUrOnK9fKQkp1K79fn9siJ+mLLeDuL+1cYWugbd
dliWY05rWnk8CRku1OByrFaDEzlu9kcSaUsXm0vknGact7WL4og4OxnISotRP/nsaXMKm2w1Tl2/
SKQbTk0jzZhkSifa+g89lp+3Hq0stmx8ie9sy8iWVBRvWXuI3mBUisohatXwfRPB/tcQ50PutrYi
Elqp6C0l3TQMhEvoZpcTuBPLhBtYWA13GCMKf+qulmvtyeAM5wPH6h4hnkFKhXfCVlcWuOD1uo/v
F7G+Z6MEBRKn1ISbeKN8G6+xFPnj5FsgtnZiSEbBVbRkmJ5DVpGpZvaea3pLa0oxkrhuzNGWET1Y
0pScNtBiXeIJiVEu/HBkgrUCqULBCcI07pwObr/6ZRgh2q4VmY5Z/hMdfjg4Q++t7R/J7TY27IHp
+fCjJeuBQTIgEanupHjWW5sdNTKgZVrD/Y5lpKQ2O4sTDofLhTBsANFCKtdfsYre5mBGwZFTSrog
ywBAggyECAmtrKtxKAiw9H/UTlgqzmCkX4K6t+KG6R4vrQXnUQARx+fZfqmip9yzJA//lY5+q9H2
ypkbRROIU7APIb12QOjMFdPWg3A4Wv/zepFnLoEQ9g6up5Ce9YI5hRPwtqbggiQsCr6ecuoEBlbW
1fIbeWQUjBD6sR/9eoltlKq0WaBYMTHUCDQMnf72btMmB/vFZkG/F5Qd4XSncBLvSjKRzfEhv3VQ
7e0TsPwMbbf/Z6w8w0GxnXFgc51xEZm8Gvv93X4cIsWfBBK7mFESQp3Ba7Mj0Cy4NWWL87n2pt4L
TyTqH6OXTas0es0nnD16dQlkb0IG6b7Jg9OLS+9J6qAGfVo0U6jJ91WjxhiXwRKY6gyrEwpiwiHO
YcCiCQZ2Cz2xEqN4+u9brLC7Rk2cdtO8s6ptT6lHZw2/j00bNDSQQBfVvyxkOZ5ThWVUIZey9jGQ
1JpBcYcLTIJ/+v+YAJcH1BjxqCFiaAM34kfPadlQn3Ni0SDtYVVH2FtS7Ol7e88b8ShZ6zFt/C+w
HcKuAOGXQM+Czum24kAHYZG0KCjEX3ndpy4OUwMyjsLi/cWH1L368hBJb1CdL5Z7uw9x6D7vct1K
/+SyOGzTqULvxti/U/L+qM6CqYYso75VXcx1Ptj9AWmEDAZ7IDxUN9ac2DPV7G5M8RWBwac+QNAi
JNr2MdCcNOhyadtpmYZkQhwTu8QIangsecqCfgOcbdLJL+8wviGawQNZG9kMRqH+cPddmHEOVyHT
8Lhm/g5sTDv5CztOT3KBNNbwzyhRGcL2vK9DcFe8AXZU/MD9KCVuesH1RF5PFbEyN0Jv6x0Fw/kb
MpsBZiMaTt+nUNy5gdEf2T5eyXdMsYIgkY2BZ3pY/C7bUFqx10DvDWiKo2OJQlMQlJE38bGsay8t
EApM65Vpj9Hghk46nlqPoo2HL083nrQWL+bmInyo5uZR/yTdGIuVShNYEDLeiWkSzucd+6Y9Miqv
spwVnKMoXquck7JeQ47EOEqTAmdwcHECFYUZSF2+cTxSb8nNCkwpIfEuh7vrQKvOZgU6DHTNoLwg
tD2n45e+aZhdtoHjB6NZVG5WkhPXW3Dw/ZSOlk0dBNW8NU3hHRaRK6gPD++v9bMJuJc4JS5od6Du
wgqq/W6LQCWuAp9WmKKNEh+Mj+6JpxaAaLv6yU4Kn/V5xQBNRyud/3ILPyEyAgrJOBPo7VIcPsWB
9hkmt03j/HIln+GQQ73ZvqEPGoMq7nVVgjH/vmoybnSvS3NQf/aJhPNmo+N+7xWCFMe7BOJbtQcw
geohFJ7b/r1Ac2rMC+6t1RNi5RSwEZdbxGWZmhj6wg96dEN7FaIdvduwBBEr9JuPKzD8G6HaYo8k
p92r8tff6UnLxiHJSFuApo05xAKm3Hj535jiuWqcwgYj1TLzRpRhWxqRpmf0VT7vHHTHG0vFADsa
s1URJvYzq8au/+YZYPP7ugunFklyzMN+8KJSaWIHF0+AaUynYlKYrj4p1UHL3oJYekmZi29ZVwkI
Q/ijcZGVCyZuAi+Cto6SZ6s6840AU26IqOMpXoRbmSwVLK+owFT0L8fE6X7iLyFB9xlQgEhP8ZY+
l4BArLXHGgV3wFaPFPX0xDtwftQ4voeIEKxtylNxyA0KWg82vBKBeY36CsluNPvquVO7ebuUAAdA
Ri1RUw2QKUmhBrNzknJhdf0Gs1xwfJfBEvF3Mk4fB+v1IvQKDzK+edb2/Aqu1FOs5SEZSRXCs0VT
Hxe3jIjfn+vG0bDdlpYsgXr5pR1yGXpfmZRVJz5Nw/biF2i3iI8hYO8Jk717KtT4Rh/Y4i482k+R
WYQyXLj6knqtaqFc63miAndHMzxNDNZqvkfdB+AUD5uAv/ca2U3/VmGUHTsrqh5+AqZmzwumiqkz
yWHQ1vIn56rxBx1YA7eh9eeGGQ8YMXaucQR/PVZK8Nm9ud2JU2ewnGEILaeXN6zu7jRWzYcX4q8k
fUxjw3H/i1jrdodU8huOSSVuCb+kTeJdL5Tv+SQWv5DcaaYU7U8j1ClPx1NhuwkF4xRergmhudGu
qZFpc1o1mpOflencSTCc9CXQV2SE2LWpE/OOq1Kgoz2kq0/r/soqeXKXBmDT/89bhMgJkasCtfcK
0H+jo8mktDKVro57m3rjyZxna94LBxfPKLLPFpdlpIiRs+V9jdx71cqRx/vgrojPfLm9bSc3zrsw
hVatZm7IPulFKuJ5R9oW+fJYaWvztqO6mvBWq9KkjS3j1eXUNR+zwDc7jKQPUas5iRiP3KFtyyTi
dhicFCkm+L9c1w6uMp9fd1YLtaUoUFb2e84AA3tr1InfbtNHqw23u6hXscT9LIGbGiENrlOQaksM
O0LbsvIlKEBbaEpwSWaDtDguWDj55QtAXAcJXCgCjN2tG8dkYz1gdfEz/mHkAlo8sQ7JdjLeGW9I
RMkvWu1N2qRJRpikrCIdg/Rv5gG2tMLoEuQit0wpYQ+bpkY7Uau37USS1+TN/RecUlSTBQjoCwK0
Y3Z0wyvJTrB4dV2KQ7cRmNYMCrtxa+tcevwcbekpM4G5DYUNs0/EbaDOWxQ3oPlX6E2DO0Uol4/s
avBJ9a8i/h6Veizy3O70jN5lt3E3t1qJ2EypBtlkGNh5VntaEU5qtNo1cKfpMTrd68mcJ3h4H/fg
LszaesDxdAFahU7O9Jurwk2B3uGKcnrmx96uiVMUG6IQrsyfX3PvwgnVLalYcuIVmVSPBUnQh3eT
uMc95FzZALAJs7k4egqRZWN+tM3esqG+MBopMsW13+AQmtpz4Nq2YqFdbsd01KiCtGECXcO8QKXO
bM0i37N+cdqAqNRk19kAzrjLnMBEjIFMW8cUmn6sNKVxvQoQ/1jKSP7HPxHIRWkbxb7noU6SDLnJ
DnnCHJ+BMLyv2EOlyPcqID6o1UOTXm34TdzZjFYXLllmchi5QCydbs7YhtcLKHpzG3dlQ9XVztxC
kYZbf9jk2O9CvNXD0eg2pQOnUtyvNMEY8id/jkAxWk0yhy928ZMAvgujjXnoKlXe4UwDJCUNWI1R
ADH/Ty7kfaSOJEGrhCVxO9wmGEz1TP7SBUT4jMrUvD8It98jtmTQ5qAh3s+C/ddbRFMdF3bOY0/8
GmOpFpl0uvk8YBbbURtjgnIl8VFQRWWvJqCk7RL6N4cDMr9+u4/y2oFqpBIA+opVmwOyo0MENbPK
ZPrISB8IuKLT8U8MOKKlsTPFF+wTXUvAvTkRbmPNa8mn1Rq5mgmrq7ol2m/xvHcEyGQIZ4F3eNs+
MJUfGTTwUAQ/uQjEL2YHFnAEkK1Krq2EpSncCoka0R5LK37P7GixUTn6DlbNZ4Sjt9ZZNWyrfmhq
vt9Y2bRqGudcj7KXqqPaKdjqcYxUPF3mvFnM/14K3VXpmYgGoMpWkvUPaUT8npJptALjCsvNbZdA
H7dvi1UYWQJ1P02aByD2tPHvChWRqZUY7WjBIOColfCZLFj/5AsFjru263RT9G1HSy13MCTo87Sv
6JIUFSQn3Yqs88QSkDhW8nPQMvQ=
`protect end_protected
