`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fzELUk1irVCjnb5/sRNq613tiOwyMNRaKCaYPZTXYpZkP9d0vEHTWFP3l1JcfSINkWA+AtN4cpkv
xuRsJ+dGYw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
EotyKCIhFyi4l3SuiXgeIutN/fnxjAiQWqBjcqngCfahUPELz7m2xFFE06ZGlGX1+9hmHmM2aiib
pqzm3Lq+KJN5YWD5BlBwlx/TEJNvuQF0ESPfVZ5DplptoWJ0+P5QAAZCLxQjbxEuimzjVEa23RBd
1zqPd3L3Ij1afxFCnOw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T+xWGOAzsDnfZDqi9lsTgiw3dfqvZlwlZ+a026rmXIXjP/VzLhA9uz9Th6+74T+5YB2CFOGOHwa1
7Xft6xm3f99T2qcx7kUKJtICvBQnlZipe0wZSLrID8uGht9j5ZVGiviMzOjb4jprpNPkdPVjRMjq
/UGnAwTnMRZs3kfg2oWL9pH+COiQZLsPR3ctuUjGjSvCWUSs7XWVy3I+rbaaKyMVXzgozc0r5L4A
VeHIXd7PGiApIiQN3zpUdVXjN6HHH4LRVsMk9uZHkRQSvTB1myIPtLGv6/yAJ3MLImg9akzAhsmF
L8C37+vfkWqG5fWaIGFuP6EvBy5Z1jVfX5nk0Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DA4nZdt1XbFiAzrWnVvqEWcCPPx5heYyoJYguRSzlzuqqFflv528w/M4xvMcNmup77g8vF2JzG6/
NgM4DL9ibaP97ozEvtSNxYGf7mBpm6OQ2+e1FkUrZTASQ3cn+lsIpuNpj9I0eKberS8NLdWHmxNb
lZ0km/4/ktAhIfMym2M=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
T25W9KPV6FVN5vj1McdrFknzMDBbw+4sK/RsyZxEGPr0tA55/X/kmD8B9FKRX//qyVXF9wtGcaSW
av7dBVsh52pbbJvdDLDWY9UvJTfAbwLNTCXFX99R73f0AJqme3nJD2qteoftiGJQPL9r4pMMrs0h
3+4fw4esn8q3GirJV5edV6J3BM2/30qIKBr5GibBd0NRZnKx86yk1Z4g606Hri441J/G161lkJtY
9dZkaBjR9Ovofs5EYhytwgWyCad+MRIQ3NaN1L4t34ZtXUoJGyvpetKwOc4CK3BXZpbxD/JJrZq6
Tqf4e0muCoEySLKPPMfTqbAmq3U0UQtaiADeFA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26576)
`protect data_block
OjfsihzoRWvRSGhUf2grJSDJnkHzRMNuIpCzmS6G2fFXO8+FYjUgqtsH/EA/U5rGGm517Qc/IxWV
NJR22K8NFpLb9/n/XjK1ZJp1TV5AcC0m5f8lyBzTUwRl+m7QTwrox67UEF+quei3YvVXAJnp06ps
40pByXXGdsTSTqTHq0X+xgfGowQsjM0D04bnwuhQmd0kM8xB/2TvUO8HAnraXdim7/Rwx3egDILk
UH3Jrkyfv3DoOtCCvHa02wRHh9OaZqiOnYm/0ylc0iu1erui2EIzUaN980I0u6glManpRj2jz0Mt
JrMJ7mKxrzzmlvfWcAqjjz8Z4KArNLSrWz8Rnz961GXtmW93bbWeNUj/a32sjHT4PU9qHL9bicND
oMPARBvGFdXfQ5r2NX5FlAS2Gpz9W7IXIIZbEwLeEQ3EG8hwJ3IrK2wzB2XUPYTCtlUT/yRp6lio
J7xfBGN4xwUakEIdiJndyKJHxBQJpJ6dVtzkT5EVVuOXQV4GsyAQOneVvwSAh3qw197W9GninHca
oX7PzOKLvs9BhAf2Pzu4ePZaHEJRa/XLP6NyLiVfEHUB2Y4xkYtuoRQxXdjI8gzLKE1DTPlkbuH3
l6eeJWuNIFXmOgr2DUiuoMHQA7k9xwXhWx6X7JNWWTIeHGKt/2YyDTv9RVT1CDCjm0Fbgg/tRQNc
4YKD/BLZIlxatvJZ/4Pbm3pUPDtLXSiqGrMqoetZT6VAeVGE2Hh4Srsz3u4I4RRWpgRZYPzQydFU
zIwYBQYWgE0DHnZd245YYWSGTMr7jUzcMzt0ilS1Y+neL9sb7b+NKzBAORsOyKAOPi3b/Ujr6yeG
k/WyTJMvNYf1KgMj3LtIvhMfTEWMBlZwj+sDYU6eWyq4Zt47U/XtvX6VolNf/E8/+w+9ysujqkfN
P6GVo2OCstM7+ydLCkBWAKFOJyuHavdjPTPb9Vj2m2eFwCm64u8Xg8PVfqr4dsA/6YVHugRjTYf2
eFgPpC2OQ/tpgdsqUWjFyo2/m6l5EV242cFdNOXVtbRXR56xp7MX0NCheXDP0cZd0X9hiN/qXMwx
CR9n6V2BkBK4e5tajIMJ2RAWZKRar5kY1B14ghQEDTrBfPpzXLZtl8mpQc3hNIILfluohkPS4c/W
KkoFvC8G+H8SitPlI2gczcUgcYlNt6Ob5XarLo/bnY9OQVF0gROR+BTqIRnsgkiZlyq8WpID2MXQ
d2eaLqtNHVus0RBQjKuPSJaeUBOcCeI8bFCvkFNN+lqB7wKB87NNusNZspW9glkCGk8CJ1eNHl4g
2J2NHJT5FPmDZN6WGujg9d/l1hTlLRVDAt6FwRofAsFm13l6HWgfXbNPIt0fCaHosEEWtYOS9Qfr
q9v+AYPp+YlH2wEPLNVV3hYwZz7rU7y3ARxBbJVb7+/rHSmCN5QcsQYccTjugErSC4qzdERY4M49
EId9BRi8taMQwC+BYVhyBoQ+yIYU1xmNfimErOFlwmTqOy+CDmEd2zIvyG8ITjUGlYc75CBRfwQk
9VBD25CCQgnR4imy+kYJwM4jsOJSaeyFtUASuxs6PLOwXTTsCvzYCkIIRzYrqMAp8fwOBctNULJ6
0qEYyx3e2WrvgP4Pv6k2yzkAsJk40NTGdm/k+oOZjt2wMVcZRrkBE8lbtGDw9b9qWidsUuvPDCnw
OPpq8Ft1ZHYepLIJrPAK4sa0TV+uAOrT1SSwERFyZRuXXUHNOi8olzIjG5hH/yxFlWGvLrUaF+54
nGl2xVk+T7zvftIh9+ohbojYVGottbT4oPy3PS1bwAClh3d41vTeUsu5Bgaa4HpZbpYDxVFxrkU4
7DLxzIvtvTUSGm7mQ6GOy6JQ+vCtnMAVZPiIiE8l/LVBoHPu6kHimdx+l+xHcXSWdu4zCsIgNTMR
8IsD451KGVlT7mnBrejnGbVtvbmyfbHW9fTX00iqfNurQRT4LnADPG2UxSabgu+Qr+BfD+wUSMOP
4pmU2AgX5UNcEbJWev0QCENTlTWJQb/g6BJM2PEvqaJYW3geD3vHAOykDgqphUcXh+CHRsCLfzqk
4cjPSTuDifEmpdTng7W4QWpyV5pn9T+7yPhL4gMYkKwF1bz9D5gRkZ2waJm3uhIVPJiqEFExLait
/Y6Skd0D4lp7tE4PWvHiO59uVfcPKpt2VR6Tf0OFTtLLhFfl4KKVlxuvN48Kt7wUKCVO/E5/Vx7p
b40EVm/aUYbUxVeE7JMlQ73BmLW43QQ2rJS6F9TinHkVwrOZ9Yt8aVn6jl/VTKSJJOBAEPDXriNz
F2ShQVfcGlWIizwTwCwUw46JuyegKYiG4f6fS3iK+MUbSTeMcODtanqPKFBiN+JCFDcV++GmoaPO
jvc/Jwe3D2wwPCfqB+ZvtUPHwmGyhqeyJPRel+ANC6WJrnuQE4x/VfsHjb5+tlPMPsUzWNtgf+Ox
VwxAPhL3nk10L7c7eokjP729d3rqNI+KenCP5URjp9cNDx6iaRSFScwZmV3eAEcK43P/cnS3lrKv
k9uvFE2j7GIuRv8PNVQuW54Z/GxTd4tZnQms7to4S1x3ajAYsO6FvjDmLkEhLi1O+8FnY/fnsy3v
TKBoXI9gh1s+pX3r+89axC2CE6kFlMiLmPr7/B7CNCr119Qqa6jftv+qhQJoJ4vFscPe69KnFKzr
Zu0w6BNkwo0WJVo9lFQYrXXatPHs8LXu5u7rhqjNCgJLOVP3OIj+M5OMTgGM3RyQQgoRk5WOfLq3
yjIJHzAob3bHtIT3pP2vz6xLYgUfkqaa2HIHRD3yToHtxLFsMxe/JzS4BsM7hzzK7NnCfqWlc9TX
Z0pIXlcihL6N7pZ1scOIvgktNtVpXHNzAq3cPVW8cXRMPWMyf2D0GiZdB3NKp5Ginmgl2vvb2pmG
aIEdlHtNWmLuu/kMolvsdZQ2SVyHumwJT4TBDLTDrmpgUFSiacav+uRopTUMms7YD3Ktq/ss79rt
y15uHyCkfs3QMdx/NwK9ksb1BFoEVpMWPap+r6KRHVs16WKc271cJ40Eu1qisevmcjYoFZToB7oK
D1KEbGEaeFhQ89Hjq0QTc79Wz71UlUHnzwlj7sEPq2sE81ef9j4VyI851KjkMoHxDStC3rwbP8tH
2+LpnswgwAVgaGXLUtHDP2KvfP0Vwk7EsJCFGUMnIak6z7R5nQoJsfzM1yjJn5WjMBIiWj2qNCpO
uY7G75VB7jo/FTUZIGlWPJvJ/1JZCQfVdmrCRDyrBvNahLUb6y4Bq7fLjPw1WAa5weIqCgdfCBWg
VPSJSiV/DaLQLV9flSW83/Qz2wacDIQhpH2O1gnTu7ECxVDwK43qMh1xUkV9neBVRloGLbRe4wI5
QWbNarlIgC9McblxF2oKB3xzlNClQhDap8AXOag8ly+vt5o/0zks2vf4SLA0kRuEkFd6CiFYl1HF
Bhnr5sHSvEd0OiM1GlDNc+sWGTqlB8RO0ibHYDrcqyNpA4PVCR1LokodQRzseWpDpM9Ni6WZROKh
NKIptJYYwyQ/Znqnz5HEDXqwcQSz2n7+ge7XbuVOWo6GqFG6UXqidUVYPJrDMxKDP1eUCbv6sMhJ
QyjCmh9ViqqHI+627SyGz1o9HEFrr0IQ+QzahjeZ/S/v6PcYmqLYBtJCrFLkX9lHyW6auBvs7YMi
Tpgpc6LBYzt8ZHnNE9xae1fT3UPEgPFwnVMiAqHdn/sZFPAeQtoCvP5IOgPl7wG7Iay0BZ83yaYt
eAXTBeH3Cr8c7dd3AC7TrI/7cWb82SKIMmZ2v99O/QQ1vWAQgHFFq48/KcO2LNhk8QpdoPbe5jLp
3W1CDeW38+Qm1VSpFJw6IFG1GV4XhoOQiw1qA3KoA5H3pLs9Q3/1sZyd8I0gMUwQr2Pn6F5nzEc8
f5HbFZoVD11Wvhz3lPOR91xW6eJeXqc+SIhV59QEVF8TD2ZjengW7qREWIRhzArpxIExuKa/LAvC
s7puOfdPxdSYMxgWGx6RCOlIaWOsNH9yrLxjOaHjcGM52kOVQ98uOr5QLoappNPg9W78cCyE8SmJ
UdSxPNOPzBXhUWuWof88TurKhKUKjO/5EsbmzMODESmqFmZtWTWowl0Al+QY9gJW55VJauxP28xq
fAwnLhX/BUAq++Hc84BFEF14IVZr2toGMbW14WClU0PwRiP+TRh14lYU+kQlCpiRWIKe/nfK2RWe
gzFrtth27p5zxmIb8bu3DvIi4t8BEWMoaS0TO0dkXxUgIw9tyzuADBnAhIEjjDP4f9UqJ2hu4Z+Y
0N/1KhMUuXZ9ELq0kRQEabbKVgSZNwKOGRMX8TwwffDNdNMBBWj7Sz1kWtXtNcxbjETO0UpVrPvw
rhc4GGMLXosyzglV1IIPTAIXzuZvlfqb7nKNvQldYYUgexldp4VNrlch0CdIAXN/lDvBjTtyU0b2
Nc9q2H73VWO0Vn8uDWlnvcqLZuTBgbY2X36tTtj2yn0UGGMODj5u/q4qninsL4m3V5aMRUX47eEw
Ltia80hRh2JW52BmFzQBKtU94jLJb4g/w6Po99OLYUGl1Nmqenhnzq9yt20C52CYYI3fABrHnMho
uS2UE16JTY/GCdl4V6PEaY4U1bNitWEhUWYg47teXmLdpkipCXvDr4I4cqYKvVI09gU0Qdd4X+He
ntjB/nIyaW4Lv6LaPHlVEJnUczWitEuU89rDmElZGXHaqD22m1uKdesr411KZI3/yN4+HXu9uJ3t
KgUM50Ey6Dpw7y+QyofGGprNFDKu1/9iAga2eZME35wizuWCTC7YZZ6MsBNpVmHv9MDAQ1RqDYZ1
5vLysoCaxZOCgR46D8CLupgZYgDTWK9gZSx27R1Ohtfn7ohCk6GG7XjAp7fBlZAqnzc4jmIh1N1l
RW6waLx4shlrs9/MNgnlDZLgKKyC0N1+lBGJMGa6tivHDq0KtY+lJTZ5RLEsXE4cxMPOo2rPYBuk
a5QkiGM91Fsafz7lP4em2f+OrSIQzc47VGDAFQm6xDuChqHva1TQ089G1jpy5oPuXOHDd91NUnef
EGWuTbLVuEx2BrhGJAcxRSCWkvPtYC8x6ORIb0Zd/Tl3vj3v6G8KsNz3YlmOgYQ1MI6YG6pdCMQz
+gd7L7X9xZYQ30RIARICsFGA3Pqn2cb93BJ0bacHgXClFIFg4cP1V4Bs9dNRequFV/aL5K6GtaZs
NgyjNaBb4lN4gY8EYxoATELFCYtGFQ2zJnjZpHWyklHSyMJl5LE/nM0pEzq2HzQ2YsiM47FvWffg
szoqxOzMCLYWZiNWr+W517Ksb72eAxRzf/cHfZ0KnYnbD0OTq2g0k5q9alEJM5M2JKSVN2BscZFZ
nNN2o7iKu3q6FK8H5M3EwzUAu8S6drwCggzXZK0EXzxiWFvKlefOm5iyaGjZ110d6vLH+/Q4BLLJ
hJg0LEUofG95bT9tPocVP8ZLxSFCF/+3ZS7Xf/ybM6AYFIFCqQ8JAio9DfmSbPwI/u9uy9s9Q+fU
d9IUkbSZCuJJ8Eoit/XIA/3dK/srwiCvXVKYgoICbCyB3AVWMfDO6qqg8x/1W9kjvbTDV+kMp7rO
YjlHwkqsL/ztfjscuD4Pledgqo8aMStgYJpINT/YaWFl4+r9nTciudZeDuA//TMTiBWhsRHVtPPc
Yl7HvM1kUqgctSxa65IOVYu7SFcToZAgoI03Xem3UX7PsuAn6bCpYaS+LEWYofWDSCVGzvQ1S5Js
dK9W3U9t9zOMKweYHSM/rzdv1ChlLaiP/fN9ChlamAHG1Cj5RSdLiX/eNTINuw2wJ4Ni8BO8CebT
UA39+VzHu6wsArVfgUVJGxcbQDT/b3wdcDIkSjLt4ybWdqQVtKiG92qWuESRdDQ+6oD/tRqHIiit
WP7lEQbZ2b+zxB8CnliKCYufubfaAfNLlF3JKbE71/AC1OFwzaTXeTgsX3DF70EnAuNULNi9i5Rx
eLeCN3Pe/3vdUQpKhCCopfRv4jW5Gd9CjJktSFEJMsLVUdJwjtL7x5vfqNZg9fIBxxuQnN25/Ko2
8GRaYXZl0XxYs/mtmylOQkpicmFEM39B242NKF2YgA6FG6Rgc8mjcE2YT5tTeGB40j56qk0RLjT0
TgT7WUxeY2aSkVp9TCLnYC46ojjgfHUSnPc3o4Mp40DVpNmI2Y82TmbHu/3RtkJyixB1wHj9RoAy
h6dsa2pxw3EcBTBy5gQtBwp1egQtM0sOvjzzB2VrqAV7Bd1ephigfssM16QefiTadBVnzU8orPBv
ohvN+q3snV52+K4rxWAWEcPFMH775pmU8UFJMPteuq70pVavmipDVm7LPI7UzTELsehVwk9erOKV
3RxKRFs2v45jHVaUSZPxtiSBXAd8YTNPkql3ayjBbl++0ZVXCpsGvMPJhqh8PMP/1fqrk2yyT34p
f0rN4iXz6Ci8WD4/Peiby7Oi8EmUZKusdu+Rh0gloXDED6GxqfqbXYTiKYYHarTBXR0LfILdaUTq
hwzfliYDk8AvNkAiLpKP4CXClkAs4rA3dZVfHrwglahJoeUTA86Lmmh2GxO/k685PMrp3nYyY14D
P724DGuZQr91GAL7qoRjKJD1OzH0deEkpJ0qEXqvrNzXU5HN+Ap1Q7nAF9ba+zb2lXfIkwyk+RhU
Pcq3+0/UrRhC95f45xEkXa7K1W41F3PPRLteOe0y9N8FhfAQv4fq11H65yoR6ENV23G6YFraMjsT
PsvDu8jqQvT7zdkHX+CIVYOcHZHjCdc9bHnFPqreDNY8Us0DN/86PWRQKEMOb7G+hGdojqeH623R
0qtDtLNu3CxaTKjRgQ3sLaTJIqVEayAkaL7wCiQOyzCNLFvpQkmtbEY7Y5jeaQ7Xzpkb0hPZGxeK
WAUqzS76Z6po++dnSn4fxfPNgAS3ObkmKB3m842xe1ruUmeoGIxUmvDrKWtERDfL9QZdFh4tk3+t
d0nyino1mdH5Zz+Tgl+xpruG595zoqydq1GMMQAeWkyJtrCPhRgPjZx7jwdUzt/eKqqU5KLtJ0gn
wiBUQFkdVS3wnFmpcib/ttjEp8roX49VDKICITjzawAwx+DfKuDG48rHDWisTd7Xo68vVdFtkvMd
bMuID+cJcD1QdNidsNdSnv7n61mUUpWZv31VTqyNDBYaA9yQBf3A8HWGHkACWUx37zSjKuD1YvZk
+YA9Kn1FfYChX1Tw8KN2SvOPlg3vLu/Gk4C5+xCxanCgPvXrhgsJmocaI9Z7PDnp5evSXX3u7dJ0
CN742ycMxrIVxSeloBSvCwLT8ecbsXEvuKgi3Iuz/wmjI6LvvakBupRHmXOmh+5h8iUX9JH4pY97
K+M7krly+NQOD/K6ik1uTQEqd6eAZPTkpIR1e+CChUuFAkqdWaWyu8PZOLPbbGJA51MNDmeG+qaz
SwsdcGdZIR/PZJksmqWGcABOsxRpY2X3Y6k3I0QRDTRNh7ODouC9zO04yU/JMSOvvoAr1dLyU7W7
O+LPa4CwYhQZSub/wiz/at8TxGQKFSGHax9voPx9sMRXTx5B70EjbBsp4+2k0yG4YrcS+bAlLdSX
kZIkLCrYm+e6Z+0f9NAlZmb0L2I7++CVY55jGLQGO5bVy0wrDvw9vEQoPDTYAV2cHal+ccP/rbdr
QstsKUwIfAWui2sKwYZYv4/gc0Rjus4Ma5sCkZIrOHZnUglo37gmwzFC7/eTh52Yqr+ScjHlKEw8
EuUhbe9hs/+FxqpF99Yf9Xu5+dYp6cG8TKAaJ1U48qfL7cIKh+GZz2Z3O6jmLYpDdlpdEd5rJkzX
BwDWxjFOJQNCH9PVimwdggW21FNE5xoDlEh5d4+Q7GM+mEPUmpqihbGc7sYTRzlM4Wm5W8g26GEy
IKXg0idbX85/m08DdIGKCnK8mJlMZAOXKMYJvoQw9vjJ1whwR5lCoaH4/ZovX91Vre9IAMPMFEOT
ibfdVI6ioKO/vGQ+IZA3psBfn5askWFMl1yMqf4TJUhl3cwv/GygZ4eAAacgCFEOdruI8WMQd3pA
/xXuCwJncGN2QR3BKEcAgu+HesHV03KSeRIJXvpeiv179e3DxGYAJzb9Z+yccinzZxM/2jYjslOn
VxtZiMRtv+yc0zNgAGSF4G01TTuEzYl7aAO/oICkmp411ATJX8YdZ2wXxG9m4QfAQ2vcTYjD/epD
Y5Hi6RHasuOc0x5ktiBPzdqzldaqqnydx06N1OUlg/hR2lYWFLc2ezL1SDg31PUP7MChCoK2DYhw
q8kA2N4kM6o0W1/wPcV2k1mAJ/+NUvWFV2WTIZW62Jz/y+rfVPuq1j8hz+8pIp/OHQ1tRJp1bSTD
TildYNrBk4X8ItMuBGCMhlKWyrsMOO1FBBRjXKPlrcYfcUoJPBlj3Ba2zsusj5RAIVpyPBUbaXWd
iWuwVev4nv/MBtQusHpo5m1dJ2xoV9cKe4CEBkvqpIbt/B19PYxS9yzJ5aUEi3eLIVkz+8us33ld
Q/YqMynzuvEPmfz8PHLH1BFE32ezBPdHK7hhSX6LHvdGC++l7Gr3yoZ5C9rIEsDRKLN72UekllSn
5S4+OidpLslcGgGH9BYlGuTU0e66tIcAs/FTewEiJ4LArIChLV/fJbSQ/fwoVa1VPGydrn20dA1M
+xzhmjl1Vod9OEEYKylA0afDcy4wYSQOixN2JekMZDMFS0ZsHck54BhaQDiJHMkpEHMgoM+i9rrN
LhTNIWAa/UqPZEgxFWQ+U1CCulCRGRtkQS9HXbzXKbns4VtRBi88UR2ZxX3fqpSSSOa4Yc1PGHwM
3n0haSMweXR1ZHU75HcqtRVUoiFFQkDcjyFcCEb1/DANoyPONCRng7/pwkqOyipi+GDgP3quAG+6
451L9qERoECUqlzu4ImU9QPYgSbNZr31I0r8cf+fJBY9mvj/6yGXSOzumRnJS7Qvf7T03DQSC57D
KuYWDU5m4+l7sziw5zurruMJ4B+kHAljfBPDrQywG5GToAAXDjcxgizvHyeC2TqpwXTyEwwuSUh5
EKHQHwoBqBOH9Sfv1VkIMMNS4si/UOjTkUQ4jJBULj0bwObHyEiIaHOCr+7Y8Gw25O3rQ0VITLE5
zREV2djInBPNqst6YeK50FqKWUJ1ct7oIcX35yZulJ5qn9wIi0sYtfAzNjzv5uNGy3nRJLfQ+d4w
3ZC40Pp6EX2FyLjF7YTNkLxfH3bcN664qwyCEHbcj+N8eqPzz0/RvJ792QxI90Ml3Wd2+e4Msw0f
i3yzghhMdNVgL6SCe98TsnyPD/gXAe5dD+Pk2QoOJUUrpW9Ynhro84kFVou9kUEA2nJW8XS13uQG
GE1KLXvm7p9EH2RMZQMCB0fzdolspXqDu16T6bwnU2Cex24zL/88pLXdNN64mv5RcEYqPZJFcUIH
H/81pY5hI95pGrR0LjyySirZG40TOrkXVd6X7BMYV2GlX9by8paKxJllfrzjqEFMyQDcAEUEQPpc
M8sO5Y9ZoseBit9tbXlB1kS8yqjdneAmcee7xUgh9EAfM5/488o/eC3w1jBM6DQj+A7xXiU20J6w
oqWScLJzbYXHJPfwlHgEwawzhpmMd1RW3wqGDJSB7fX/FyhrraOM7zCmZMCIFyx8vovVHd6f71R1
Ld01OnXyEvAZ9MAedoOzKyRDdmOiylk2oBOLwVz13CB44o6WKZW8pbJNAO6L7gdoZcsvoY3FDHyc
s0rzJuZovnMq5TTMEbtMACkWFxeyiEMkqhHYhqg+YB9vA5uAUODIAq9tpg6fbRhGNIIBfHm2DtCq
vQjdRDGz9gWbOf1BEQzeFm/K/oX90I8YFJiyrcoolnUTsj6bqCaYXRNWegYdo2aRfyPIIIfvWmAM
U5S9H6C1FBt7gu8HrmwzdX7RBWLEX6TNyC0fKs2ABqcXmetgDjzCaYSwFFmCYIhurlDTMND0ZGIO
yxb1U5rzAIOy5QiOMNUyTI88oEKdtQnofocjMWB2T4kerCXTSBzyNUOT2HEWBf2c6ZuVGuS1KJF+
oYk0m2VOEsxY34B3N/cSD9NFfSXpT50WxLDsbVp6K5BGiMNO5uO4f1l28C/LYitiYBQTfjXv4MnB
xAOzGC7d19R2qR3cQ/MHr3y/DSxEdAOduuSNEwxDTtPEvf3/XK/a92mNOuSINnt1k+bqBFoEHnXp
pt4lnM98CBmxbgHaazG+2jZGC+BqZUFgs76bQ9S9Nmwg6qCw+D3cdahJcN7QaTISct9BXI2+zpWy
JhnYax2+BDN2ImJQEymmhXuIsteU7fWJaoqMMGqZO2BZ5qX3zeQKn+nqVCyo1V2c7uy4l/FSDvMx
wqdX1BIJD/g+L6K+3Rj9a98UHg9JecaFYaDtUFFzhatSPD8lVTdfUgInBZamcGTDm265O+8kDbsB
VIGsjpFCmHgdTjtPmUzcJJHbH7qif02AFTRHOy/YxZs6Cr3ulVV4bxF9G1AX1NIG2e9WfEg7KB5Y
4NR51cpnj3fbMpb+eBT0O4STguzEbnj8RFSAZNeNlMJDMk/Pyxn4+Z2xge29nXpdbVeOd8z9wwHQ
ZLEHBIsML+VHT7picdvq6EsvJMMF75dwmrXQFP7UvEN4KZBt5hzwiinvy1bkYwj1pl+S+mI3UHUK
0hFuS/vli6iBMyiNpcus3QmOu3AlVUXYbsN7ZEqQOhjVcD7zpWOnzNEcCgOq6iv3EOE+5whQWEWt
mgo8QeQYsriAMoYiHT49+JfXCf08Z5Tq5+hKgXe5qJcbj38zg3xvGG5N7pLTHeSmAbbYOmwwI0Jj
wVlO13EJHmktASWtnfB9E8f+nTEVb2pmNON7eJsLmMYronTDVw4HlglLrrlaKsbjqjvGpeLWlWWB
HhGXsip9zxIy59c/x5dmPKV7n4Z7+00xn1XjUD4Mb6x2rY3bI88kYpjEV9wkw2SyjIg5c8H9CzTo
xnQctdEohO1JBRHDmYYakeMOgDTPW/Qvp8beaytbGq9w/B7fcO9xifbh31SZ+cXedeI4Svw30PsB
Aflft3kL4D1zRDLRSblVxldbvQspjUAizrEOu6KmEgAvg87TxBKRH7ZXCnsmIODGHgnInVp8ncgq
hPwTnIF0LTf9NWFunhYpQ+vVkHbXojCsuo+/mK31Pic1QZvtmZ88V0bFfa0Mi1NVyw5Z2odo3rO4
lzYPN+EaHpgw7IKIoik2Qyeji6ikU9RuLjGfnbXm2aVOmEBCtbF4U0Em0q97Fk13fxk4JHG9BJdS
8Ht/8up3eIjCBHWbp+16Eg+IMUjN+Ci+BcpLkgoAMHqU1xLqZ5uE0Wmpqg1TnkQuw2UZKWK+IVoZ
X13ISjULuPgR7zdGo2CqtlvQ4emT/nKbDEoieskE87l/XbsaiTmbxGhhg/HxxC/68LDIgpnVgKZP
ZYt/UAxZE6ER8GfDpB7MWBMP9QDXvNIVPxJWHEAtGdbDtElFyh+mE5/tiXfMdH+lpOOMd/AuFWB1
VBgsGVZlzfxkkey9Lg2tmEM8hVzZ/LCGmdf0VWXeExvthwW3QtU44r7DFN2p18YALCjC8s/2mdDa
wjzL2D+Yr7thxPTa9XMbFquvENUFTeQue3Iph6Hg0ehQpGa8vd+qR6Dy6xao/x6EWbH3NxW2NIuy
+lkLMw/Jl01YmN7LyJW/cVXv7PmgEaXUpJIEvLRkvVuP3igYc7PFuham9pk8KW6RnouHsyxTh69h
949RZ1iqsHJ3uptfOeMBtKOLcoBJLRgkmphjgNelzPI0CEAJJzuRxrmN4dBmIEiNwZ2X3MNTjLBF
pii4f636H/CD7lYKsyCCxpI2kisaP1BTDQXyzsbhT25oekI98NE9SQiJUX4M7dHcnJxsUYkZtEBD
ebU1QC6Gmws4fvcPnnasJVKH6BbPNjM1t+ISE0DYFtqitmiwBHY80ttCYvQxw6PGMrPpr0s4B4PV
sW3/QfcBIAsV/wBAjCqigu/BZG5og4FqbYmSr2AIM/dmmZ9ywQLws5zS4eLD6fCQWdIljngB7Vd0
hzmCzxYZLaPfyV6sv1ROV2krpPnGC4/KYQ7zNZ3yWwtPTDlB+a5qz45meFHTUDAUP+m6jSsJ8UFf
F8LNgDkeRt+Iq5EBO1nRmh5xaS3b6TiRCNWVP15G6El4Op9hu4+Swtrk0VMluTu3e4mGaZqRcXMq
nPuH/3YUxJZj+uN8eRDJIBvNqcIL7WcK88keB4Nm+2YUhW8E/9aWPDR44r9OpJ0UJMLb2MK8QY+S
tG40Y8n0CtrGwZsauVDO7jAoGq4MUjmX3ZqeuOuieUnWesIwruJO0yBtYL5JOzBFcyiCSpcFWiRh
1mTU+pPO33fb9NtRhB5rLe9D758bCE871EZNe3eqTm/DlRn9zvXf106amuD412v4cBwU6KPeucvq
Z14zU1RRgUnhc8lw5NHaf44YjoI2VeZg8md2QC8vpFa4qBdWOQgx15++AtAXAJzK+MbwMXMNZedL
UWcrbdlQinHmSknqSNxAbk85ggVLQ3lA6Q9nvTDoyWrIW8M2AcsG8knDAFzxnukCgksPPadoTiFA
fERlJLcoXTMaG+F239cyrQdDhxdBR/mr14+TdbQxcNP8+/KimYgK8XtwbmbZ0+34k6gTpx5xZVxL
M/fMDkLNk7KcTRm/c1XCZNaPCPWgE2So7/AnFsSeiv9J3tWigZxFqkTbP+hof6R+XDpQmSp1hZ0G
OcM1i9s/JO/3j+EOeSDsTewpizw0Wc/FbvXNE7lL0F/KMWvlKy+BSlc0sevepH/BgMDJv3ZNDHwp
cE3VW3DzUNZ2ADgdW/iMI4fNydYWnLyhGlk1b85lV24OcIRUGSe/3Z2cZlTQ9JBjj1G4O5WKuY9q
Hv4elg1KBvWVsd3RoMeJiUjBpJTzd3zYFLvbre5QsG+oKxHJbuo+pvn1PyUIn3+6vj+ObcZYd8JM
NOP+jRzcaDJTJOBiVI67g+hDggAc4WbjE5JjfeSfg2PPyB0qjObGvznjE0CUhFRO6A/VpaV+dqCv
kyXQDsKQqslj3ybf2UGCmpRuHmvFFC0SAnBsEVHZeS4WHrC/JIN3y2CqaENp7OF1ntZIggae6pcF
Un1utav0bcpvQYwDNO6HZZn0TlieL986/9m+N39+ko3dUt3kKhQ4yG8tzrcj2taEKrsF5wX22USK
mND3nbYq/HQWQvz3tbwZFqAnNHIuC0kyy3GOIQzrYJWj66NDB58atX5kQL3EjYglqjhM84DsnIQo
uacpKvAk1cxU3ZLOf4ceZvgQXPAGiwSleSeuOlSXMxEfafNAVILvDGTKXGNA0SCWd1N9YcYWZ66l
EW1Kr29g8h67ioBxDdCiqUDgZiXBvXuqOWQd8u2kxRO6CinFYZMVOpgDvTw4cBtXyfHr6UvMBuFI
pi3mzuwlzuwZNNQUHAK2jTUsNUOwycBEXWncCFzUwIAMww+CPY98aMlge/8KtwaH7obR7rfPQIVy
fyZBQmuNX+spmsirQOBZlPQtEId2KgLJM/p8VhfZPz0P7iu9qybns6QQkZLISB4fVAK1DCOzpkpw
U6TG/m6N6bePRdnLaJFLhsDLTHu/yQdPfu5gc8ACU+TBDXp6Iku0cmINd6wgMnOZMFE8uu2AYMDc
eyn1ObbNZw93+Pxvs9Pec0A1+h0qoUUuknW4mVnkR6faFYzXwAB0UrUp94PI3dYNAFkvttfwza5B
dm4MOHvWnty2P73/oXkdlbuDEkU2w4gY8hFM/gOD/Ucaxif4JlURrJP7ZNE3s3EuU7eye9wW4WKl
d/elfdJxWcDslkehlAq6S4xkpJ9stXjuo9T3gjxlnnNgu4lcOrTfsw+gXh/tDxcdAGkh7nBTktwD
yPZ4/fKYZUNouihc0O3cISC9umCH/IuubTvKDY4SfKeMwVNnynl27UvzwrAavln7DzdUrD3AbEd3
c8R1pbmc+NxSHwDUZf38OudRj0TQS4cIEmOOFpLB2br7KDNUzCmkY1CwxYfY7YbNQub1SxxSAEg6
CeqklqBhjRIu+uIrLs9hxMkqmm65sEfFAvGav2uMAdRdoJgzLqONbE2kPJzQxQWrBdAjajjB/aEx
3RKshSFcqJMgWLc2XRZmG981uhrw+Xy1M4yYPi3mp2LEL0YiaSnBcGwx3QMSiYYJBbx55VewnkAT
foJ1XfTL8SWk9iP2U72A5KOmpkrujWUOdYug9PDDdGdmgvDha+bHqbtlCoczsrSN9F2g/QQGzO21
sJPnZNx9imWVl+oy3BAst6iy4gzYnpYvZK6C7OrR/yayiI59+q5ZOrj0Wgk0WXxmRbqakYfOY3lv
gzE1p1iYuyXseDW9FkdET4gD5Rgf9G6EDPE5GHGNj8VyGlfD+yY6dZIZImJmO6bqH82rfZfuC5ig
+SR3Tho1DkSog1yRc/HwYrGQEwVYzom8UX6LDqZjl9h1MY8znGxIzaZ4bkfa4sBW6r+yeY9yClLS
ukzefOr+DQKXRxt14+jb9g0/Dr7x4K2q65qE9MzELZwn3yZklvHskShVqj0RK//8e/pBr5IjWQ0z
VtKuGyA1wTOkI+t+m2u9maeb/rXFLWPk/9lbyqyDK+AKHVPDcYVu+CaG5+orXdmfhyx6c7lmTcZF
mdNNdic/DM9Gf86unfnc+JRS+ZvMBktvBTBdlqxZ0VtAt5dqOBiiRCIurHRkmnqm/iGUeaEZwGJv
WAc0UYklG9r2ALzgs9lZq0sWzPAdVKWPdo86ViG2dD6/mIWmTxRO+Oy/iC0eoItWGD7o7m0nGuRM
Z0TI1iD14G8KWMQ1q+7Nc57IzP93/o1Zlf2R1vQFWIZwvOr3GxwMDAeJBHA0XGKUuGlLQBDJsSke
RqmN0gdHD6en5pgM/wkaQTwd/qpPH/A00SnXeHU8eLwG8H5+HbgyYIfDz+CRtmWxixKjspz9UHRr
R6XzUK6D8OzpRubSV6q/KdlUPp5qCYzFTExyiK2WkncW6SA0Tn6POHMn+6SeDT6vVm3Zx6IR78X8
V+DZbNRmxNQZEnMWom8AbgsMXBayQ2Ammnae0VeItp51ibT8PUgIt/2+fHq1fJtqdmN8CY6qAQKt
394b9Eup91LGX+TSBBrUwCZwg5SoL/zRcPM9c8KO4vkziu2n8BZIdDdLLsGNMx6QhJLlZBMDaqz8
ZW7SZxplaJdI0gmlL0IT1Nid863sd7N1CMvXDHiFfqV3Nz081LMxQh/1goqpDVbEkHPLgUaHci22
G3ykAVb7EpvZhNqswDvOgBdpJJF9qhIsN5f3r+7LeM40o9Vn+vEa7ALIwZpJCUKQ08I4Bj8mwOXX
ZCdtdrG3XwaEf6+k2H0U3hfckItrO2wO39sa9C4FgZksgPoLBLsBK9cICL0skO7En7umks5ztNpr
lFI3DbU9hBOG404DtD6wbBXFB7FfNdnvt4unpsYAKQ/jkileN7ohboIuCCntM2W9BxuhDgwqMCvF
Bv2sa99BKi0q4Zp36d6DPvEAimMynYizC+8V+xKnkfct+lYtlHMZKLkwazOSYusYMoeZu1h2Ylx1
0jwqdifeuhO6htIVlVVH0satQgmLTo9y5D6lpAS4yjWur0MlIwWgIX8hPZy3HboBHyLfpklXJKll
qLOE5f8kKZ7Z8Ri/qnJDgYVeFkrho2nsy3AXdNs9uq1xHpZXdGkVkWf7TsKFCwS44J48Nf+ZVhZ7
ZF0CeeQewZG6a8eOhdke79YFzCGX8KQ8tFlXV18o8jf0L2w2kRwQKCyAWKuFXv9be/vf82Y0EyL7
VA0m4C69JDu/+4SukV2RCd9I4fZwggetbitUI6czihM7RsaYZ6yO6Zo10pmYvRxPXxnkNP6IwQTZ
h0vzxaLxx247v+vXvbbgKk7c8fPwrcb+7a7uxu9Mx+5o3yAtqV9gKMUQuCtOjicDa8jHz+0yVl0t
nbNpuPRhVLprrUrBKEX01TAsbyxMrWGKti2ECqpR7hmWW3ZnFlzai3Lbm16ivPwJKIiVB94QOtud
HyTeHOlxnKq3U6MibnWP05zxeZ1Dzue0cDWsUD1H2DHx6vkdYj9KBzDqSUqr8XOGySQ17NrUNcBJ
vIU4TsUxp8dLy7tktiYIr/G8iFpp/6CaZVZvHyn74Pve5juNVxO1e0Bt0bG+yph5STgl8py+/vPc
G9EX61Q6w+Yj21kEHKMaYk10r3Lv0e/1/LxEusZkeCdgBmWWGJtA/+VH+n0R7bkvHihe7UfmP+dd
aYUvw/N4VnMhL1kaPnA/e713sJUUmEOcjkBJtYvZIrLpMNF6X7VZdZyFSj5C4ZbopbhAHZV7sFl+
Gf9OhCE1w3xcqvP7q8c9HMRxG6dZUcf6xqvfc4Vb64Fxb9AHj6T5MQY2jx2XL7GykmUVPuy73LGe
KhhkNK1hOQ208Ztv/J6FW9DYVQQflyGewspMAOanAk/MttbZ9qee5lp0UV+ZBFfby7ah+MDSOf0M
rPAYzp54L/aymH47kSZrpTyTxbRRvWwGK95jHhs63XAwGr3cUpaWw1/DfD+h7BiiGm0NpfmRMbBZ
mzVcOPDqBnhltf7+D8THLNwWyLtfWMYWRkYQ+zRHxkDZiRmXMiuyuQ241dcnf0ydrcrF2MzF8CX6
CZDzDrDs+HpLpwlU9+u3/1uiYTSdc3dn+mCrOljRiHyTHkgDq/vGRyiVQ+fmtNosGzzBFsOmouFH
ouj/y/5PjZ1V5Fmq3uez1fVy/Rb3vUBY4RRUKsIl1QJ43Y16LyP9N/VHvXZ/jI37oGsLCh1QhDHQ
GlxPRtoZCe0SvQmTD5X5JAPd7RZtRKWPCb8HTLhBWB6XProRzG4xNpC3vVPLG2T87gnIfM2ETk9g
31frbEubNQ3UG7P4d1RRgAqIChc95c8b32id1PhVJTMIsB/+qgeYAYbdpYr360Xn3n8TDekpBZdm
Z84S9nDazMIe1MMk3gfmV1AscZt20bFtHmGs89ekVckyuxdLMg8hc6PjEUThQUsM5Wzty+Yamhiy
B31Nphdk15t5tvPBoQ9btzVs9cXzAyCfsSkkzS7cWPWnvt2m/xmHYuJHdWKTzLWljBP4irptDhaT
2xQYnYMlagQYa+RsxrUFDLaD+FtQz2l+kO/rKyBcYG/FHkcQ9d9kMOWV+Q0JbBfxKEGz8ZiVCbI0
KljEA7c5kJM1YmirN/iX3rIzEgFif2nGF2C188ffdvrtGpFz9gz8ylNdZrhDZvRLt8S1s6Dw3pnr
RdQs9g2XB4XHIO+oVQ0iMcSkun/1fBov0IC5XB8sESStTMo6ywYAAhASuplGmfnUxZRLmV6ktjp9
gND6XUz1XsnHN8LIwGC++pLSHYWHoVlPqJdZTfE3a/5xXNyYaltj7gZ1WYtncjQDJemFoGonxFAH
dhCLVGMLxsj6XuV+UHWI0ZWjFJq1XoWlcWFKEa4Dhp9Em73vOB4E7x80WowmAv3LQ9j0W5eXEaK4
57h3QihUwGlCIF7dQfkr6bpUhKE8aE4ClwL3N56BxEC/zvjtXEJ3rCx1TFCu2fm+NuYRnWDsIXv7
x16cm009vkmylE1dPkczC/ewItTYY/ncrhC+jeK3dbT4fvJb/W6uSEOTpve5qnVTXQKeKygSIjBq
X9XQ9S9MNNYsQy/mAEBiorWgtdvwSFnhyKL6dZdS00pZXOiWtqI1rKWZ9mKEfdXDqGvbP+UIU3tY
AO0eMQdS+cqSWDZxGzf9wMnSyavdFxiideOsvwwqI4/jpDuX2X9Nfj9h6HcrLMcm/sA+1iE6RmKu
AcNLGUUfvsR53SOZJ3ugHAOHWH2/NoeuAy6Deue5DY+2Xh5Yk0a4MHPpQoKTo1io7PVQz50bxesI
WsD0ETLytHrGEJMPEeIiF/6f3LchXW3WuUtvCwKL732bEGwNph6PP1AM4+gQMyOjirPa/dpiI5tv
/Hmx8C47EBCeQigkJ8K6KPLSFko9wclF4WG/6BW0z2j4V/9DqJFPRKp2vPPauWG21RzevYNu7lKZ
WuLUQe+4K1T6TT4CWW+lqb/BRN18jqswe1R+UTxwqJNiJKQcI/0ET0vT6+ownNFv183V3EPeLe3o
usSbUT63uyD7fCJvlwR/qV4/0XelEw8+KPBlS1X1YCVUd/526hLN/5jQ7t67i6XxE3runIB0Ic3A
bpaGNGmfZnn9P9H4Svid9eqJeW00B2+gAqCOW/h2301iQN4GRE1R6e4vBiHIm+GzSvLwxvkRfxlz
5iyVQDPCYUEIAFmceCgn1EuGJxzbMKIyhtiKOVd+mLvY0no71WF/8R+CUpbA9PJ2Od/OxXhZCcF9
uMONC+lT+dRNDD0IbTp5mXFWV5/USRo/CDRMaB2krngD7AJXPO206+9jlpWb4BzN2L2sYo/BTEPs
BmSAArfI1xeFgi6rXj9TqKQ5EvyZTkoPdPiCtoaPZ+KzJxHHT+99pWIOOFI/NI1k4crN/3laoNKs
pu9uFuEK9T2J5FyloTJHCKVjBOjSBCQujKCpLVWGN1KgZ+PES3O9Gwc0cjhVadrN9aXvJYm/xoep
JEtYNEwshyKsZ9Yvyux0n954iX6ID19T0W+2Hr/Ke2xt+ta4mmCofMW4hnAcXvbyVGkDXv02LwnI
UVcAwkfpPM4Dv4QluvGh7mNn3WLcvO/vs7SipgQ9pZye92TsxWeG1FTgzcKApkNHdz20PlmO8cN1
bW/sMKAqKbUkIrXKN5uNj1KhpiwopaWOMsse02imlkPMSd6sH/TOcnnDar0zS1gz3bs569B9Otvv
OEBppGPPbN1FRSBnzDVZTHh3uCUKsX6y/3vKbZuitNq65ozyNfKseXaO8xvYvu7Ur8ohUmb46kJn
Z21fB+3fdczNaX6RoqNYBOnH/r6tqcbXK1U70uLiYW8TAtPyBOVpmlvuqiXow/ot3y/JY9tx/rjj
CPNUNjU4krWcU3w+rl1HNBJtIzkscxnLFaDtCCzhfAfsbDJil0900cN5CfC3xJtIJHciWcdHbs1f
2/45on9iR9GuLNhaO4eBrX7r1hN96ElRf+k0eP6AFbwX1a/w/RjLppgMlI356wfykszur1Gu8LxR
xhZ0hBlUauC3pemzJQvvaM9mhiZX8bA1Bj05yqcm4hdSV3WU8xlcFop/qQZy01TgVGgtiu0hoxqJ
rFrC0zmnRmlrToJZPnleCaUv/uhcnbd7ujld8XyM2UQs86KyVQ7krKp+KeljNPUjJn4RewKph6PH
s/0ELpcrHx+94Xjn0O1zh25/BWYDrwhdq0XAUIpyMbRN2VgSJP7o7L8JWrvheX3WKm7IarEUasT8
bZQQydXQ4m561sDsVCeknC2O+t3/p/Re4xuTVpZ+SP/f/n9X7j/KBtYM2LX/dvewpKx5QEFSwAUz
/1rsi2fpldx1Y063UFwyljXLipOZ53kdq/dC9g4ieh9+95z658IVSpIB1k/fzzCroE7ZqKoActL7
3Z0LyeCN/gxyUDo05n+d9zjrvjXK0YaXmHamBXHNU53EQKX0P5Yv8GYrvzAc+2x9Krz02K4X3O3D
MWzyMSK1oyElpQUmLz7sT1ftQTFn6nctq/0LfDSnH7/AFa9YE03Xi+Q0ZaEgCHTpKsioySzUM1r6
t1856OIwGQA0S9PbFzkPoaTxqR97MbiTJTB0X2kUD1485N3HKPJbMKRerP8MV7qoZlBH1eQ+2LH0
05oMO3X+BXQZrcuN8pbdirs7LFDNlTUfKKAe3O7vyzGKb9iGps4FRWnj9TBXHRJsYlWe5qd1tmHn
fQbrWQX59nIChF0vLagVr2QnqtQMR7Ql3InBG9OhOGAqEUYG9oXtRQqpzYK9NY3wuong1zdqT/PY
GRlBVy4gGi4XtbxfyJCDQC20gHAa82WKJ1wy/ECGaklmhFCicECTHvPgJtj6h07VAfIEF9HEv5yh
4V2/Y19MqhEU9OzpTR5IZPZnlJUGPB6NigX6OM2DjVMbIzHi261aoKBfLuokSBez37XWKpe/uwJ3
jenf1wuGlBqBk0Jvb5EjJMrGyAYTEJNFlWGu7Ek0f85FUNgxfHuD3A9+ha8/e4Ve6FsmjvjhDp3E
b67i9cTo4KacnBOgH/aV3jt5hqG7DGXyHYzvs6icuaV2jhDXuMWGHxiEc/uImDmctMXA67vOEa6e
MoB0MxClHSDnLAGMLuPqqFCl4DJxn1q0ZCW4CWAJMStzxWaiOIkKTnIGTCfa/kJ5lWTkLr6c5GiW
vVZaJHfae5v8GZL5gn36a1TsmjNJJTTtt6zUwN3PHT+yX2ujRzCF6mPaS6RsX2OcqROhMQ8QLWnf
mo3/q/AXKGWanb9bN5X+6rOX+8t9TPFVZBarZv6rHnAfYP0WYmw2BcBz/9ZakH8OSsEC8vRMjnD3
32vw7BIaNfe/rrr+RENyJ/jo02dSjrSMyRQI1A9ADyXAfVjdCQLdYLOy/X02/7zZeraB1k28v7nR
6vTdCVrC+5ceSOpZkE57FAuT0ARBGFsbvBU6QtVYHPki1iQn8r7rIR62aWZMKeADA+1cOW0Njjg+
YV4+jp8Z8xJUsaUve3wPwv1hEqK9n54hCRWV5zZsqmk6qIZrNvdWMZseaF5PkZYBm5clNlp+LUbw
iPAMpx35fqNA5Z2NXHgO00F4GtHZI1XdeIbSrFRPLPQqFeaJKTIygHE4b2b2WVT/Gk5HENiqJyl0
eeS14sNKR8OgkVjG/e4XvnjSMI+ppLZhR+sIr5nQkaVozwcL0MS+GJuinOs1q6JueHD8N/Uwsh7t
5iy+aLmkmvHeyoWsLduw/yZcdTnsbtdsPIdWfzpopoegSQmDfoTN3xBc5qYcIxyMjpi2Z2fjUIA+
i1EFW75B++58iriwM4BJrJFhZljdh8PpnFUWx1+JgFqwIClqHGNt+S6MWH6bMpko94jp3oJUgtIb
YNb2a7EGvyx1ELIxKtDJXUrHhipZTnchk/357rkrsENMZ4aGlG2L4B4/bVrtxFMtu6Hfa/8+k4Jg
ltFMivyWkEU0uWd2y2f31KWv6Irku7TUk00HIgpM5WIwPgU3NDGX5Z/znnvVVKmXenCI+UE6AVOA
m4NRDhx3jWUATZiQTeksAdZBDQivl21CAjbHgFnac/gl5xfKBZgtazeYYzF9ZEJlNWNUPe26CNTk
oaj8sBf6dIp73kuONniPkLH0Mi+3pOGUC9uLG9QotrEHYkozdXXQHJl05xIHzrlbIxGjTcnTex3s
qwYzCYk2zYaKIoDCJM9CBJ2eKj19q4zvAbGSBd6Wu892dkglTiI4/pG+JwLwxg5t5gx3EImhHXsF
FZKS0M3a3Q0Wfi8bYOW8+S2qOcRwZ7XNGkMpURK9qJTQSOWhRanBDGrtAFGQoszGfyl8aYPyfoQW
vuWfzgmgyOI0TQANoBboS0N2W9gfXPKvKfBGrreEfLHHCqMwI49erHICV5WklhC2pA1t2Cv4nTXx
/2nN6WYkOuYnTJktVCqqtM8OQ22/dLdCVBeJe069Co30o4Bc0opTevRdXsXu1laJyhbawYjKfu9Q
QaZrnI67+1yJ4RxhyBW8YgYSc8kh9i0Q8AhF9P3k+O1W3SeoXlKzwrTt1ok/4AaffNfBxtkZPeKU
eexixinMTVlR0BY2cjeJm45GbpCAwrb1gUipBgROak/HcZaM/Z8AcNrDz4eS8UBl5qvYRasnsX4O
aVOYYM/sHPiwL3lLLEUVA2E7aRtYhHObGploid0mZ8poQ13ghhuvVeU01yoDRMTTSknQJndR0FEz
q07yEDCOOfURDg5OU4HmIUpVtXDqeDWM5s3dvgGix+9C/LHLyNpYh4HXwJ1j18UZwe7Z/Jc0FfqN
OH1B0bZ4zNakzPEQJHEFLu61IXcFsT7fkk4fambbqprtVlONUrAcvvxcEOb+vmuVItSH3zorou1s
vffF/UAre5sSo1LsL+9UvNK02N/xE2oQIdOvdiUn7YLhXz2yUvZtkjAxsHh6+6DvWgv44U4QOYnA
riCshGow6G+32ayym48Jh6m7j++eWHDV0Js+mknQbLZ5Z62826vv5eb+ckn8aSBuCCGJkd048+cc
Z3Fvq+RpF8myfUle1O4FEjrgKrOYYcqCQHX9hY4YM1V7mklfJ9P8BxKm0AKFSN+oHx2r+hTHygcC
KPxXxCz+z8Jmp/BYDbTMmrvKeTNGM07nfLtS8bmvFjShYrH5cjKgsjgQxon0JM0YCYExVEBZ/eyz
5ggevfSTawZ7fztNjIqPpCFEKsG7uPAjqYEdrb20iFANH2qzgjwBYkkQElPwQqqbo2WiJJR5xu8g
4WlpZtjqAxXacMEKb9DoQEn4nWPzxSPez8t9oeNODqW+LL9u3QkacVJCklUQ7NCwWVezRbZOAon9
VKQSZoqfJrUgaO4DRxG0CMUvNpHl5TitbKUp6GepTCI5yd8Wz/S0eIyeVYBwlnK3e8fI/q8MBqmC
yFy3WWsDAxQ8YHaXLMS5FF/m7Qu1jinBytvXMWrTCF3ZYUwd4jpqu85iqv1/nDhPm40hUcxPDNWY
WcQzCDGTJiyez6yjsXKiDyJJGW+jHeH/BEsbvX4A1bqlsJra0UkZOC4MWlhEjBUOvbUHjioyF6XY
Dnj62CDRXmtPQFbwPTn75SM1HYvoBefgG4LPmcUCiWvS5R9vLGzs+80x15bOWG8i5hwl+NP0wUHo
eGru4OfrkbjuP6aX31bavy4iSb7oFHlT9VtcL+GvFGbLNImRr9cKz/r0dTVeBs4rXBEFvKU/NyyK
+miSfdUwgwf2YG/wF3q7+zEwA6kHsjYSxsYaMPswjA+VDB5OAASu9uSILhdFGnJ34N9jpSUdLJI7
OTGtNx+8g9v+V5IGIJ66AAFyg8WsaWmOXjbtaP0fJCZuToqYm5mzevycNcbXRgjIVDI8scH1b7pm
JBibe3f6TeTkX2NhBkvnTSEkkG1mZZCcNyhRzk6EBgaJyEZ58YbmplW4pD3aK5c1uOW5dhmb2nuf
F7MRKIeHnk7EAxpAkyYrfCmCuAPmITRA7TIwVJwZ1DP7xdQoG9fGdJMM9JvDLmyWFn+xYMBXwULh
tRF+vrn+tX97BtjXL8R/wZ2f783NOq+Yi0HCPxWhV8GWz4pGCa+GV9p4kn8Rsx0NWP41VdmNOm2g
/WOu4E9MOJN9p6ZhPS0EtlSAVDbFGWOfjchjnOb6bxz23xlBCOWv7DJfATHtC4hcG0ZUxQWcG/KP
mnFj52AwTpzEN/HeRr0SBTj/dO/PzEczU+G8IGYxVIaDlTHhhTw6RHRiNgDSJsSZsr6tO5Niq8CU
kL5ZK5vSB0/+R+0IneQ5NOtO876bK+ZCAZT+IaUvezbC9HxhEjsJ4p6eFtwh71x1VgTIgzcMz1WR
6YL7h5MaMLArdACUEste+2zSS535pcYn2XHqTvwHIPJB/Jn/GOV8wEVYJKWXMqJ8y5+42XJwjK5L
6EVdlTrUAf2kHJJFxW2rAUTqsdf7IttQEr7OyBgt4A8rRDD8INh+uCClJy3U3afP+/WDRFEMYyNl
D4/vqbr9GT/+9dNwt+3XmuVgPiucLsJI0iwYqvGeqhWIgsbYSs2DPe2gTBuR/9VpJXFhcadmdRIQ
qRZN76YHDjm7tlMOweGHGHImLENWAvOphP+/jd11T9UdUtYNFlgmtKoNo0wuxOziVUHfEBAKrNz/
mHnigYcqbyTx0b1D4a2mjvdQm5EyJBVeAqGSrrg+luK/bH3IBv3F+cCnxqLZ1aQGFWmFtWnEBB3i
d1M4aFsGmQiGZiGkJ/CFV4y65jy/6BkvWQ/TSoJo9WKzsjeZUZTj4wB1CgN2QL9+FMopS9XRKAV2
t52jq4piFWH81aMUUxiwlK9VFuCXLxueZno1N2uIMeFc48YvcbreGuzoLjQtUU2tQJPKgm9uwioB
KceWdZD1Tgcrfz0Laq1ri8YEfUhawMXnxbwCkmBI0qGGWXJSdz9ani4Ujebszelje49Y8G4GxL4l
tArnAMtyYKfS7UFZoVq7mXKC2WrUSsZ98qOxMv4+BcBimA5lzMvkX79mXPlBgWvM65FhHtqZ4VK9
e5gQhXSNLMB7NaYEOQx2pQ8ciyUlYzRlc1GP9KqEQlt8WvYYh3Lap8TOP9bDT0iCBwf8nryRjn7+
mo6KaNMBdGEyrQjyPfTdEeX3jIKCVz25W5RIFzNjjbMvQaNvFqEpV33hpeWURRV/IBMJghHk+3cH
8xgHpgNlqim0lj9pCiJkJpCpxRPQ3klUBgJNUr4vX5GD1ewVI1CYpLNmzXurAwP/AXVzwGfDJUbU
oC4qV4c1DqybNrN/DfJWae8ZEJ3txwhMr3ZavT75aZ45ck7S6SgTErfBkTIWYocY1VZr3cpshSFg
vli/tWynYDNIPIMuVuZ0mbutzZoQHbeGgmXVYWfYz9DCBkbaimGmrqvhTxxIoFoFSN3Wtkj/rnzc
/BTBR23Y8doRwLC7BbI8COzLXMIBtTpsMAa/cPm599AuTjlL89Xwr1Z5Hu11j1eD+vzW7NZDFlX7
1ySD5WZ3hpS3k8X+g5x3OXYz7hEFtrAvw+HhuL7BDLrpzVia2GR/0+yuNW3FhlgMF9ymG0191Ylx
d9uti/okUWiDJpLQdOrtXjuwyrzqgyHnuV7VjpfqsDhz6RsjmMR+5qdMNIJ89pIGvKb/DxqUu1iG
AaDR9tOQMN0dVqgx9EIUwpLFYtu0PIBAZAgiZGwDb0YEYr1DOa8fJPoqtvCIs+pQqBDN3NOfiCGi
r4YZOCbR2GQZ69YFSJVRVUtWdDVLQw4TPYE2i+0pZBjdAjk1QrHs3zwsowlPgA5tImsgiHTW7ITJ
OJi2a27ibsDR14Lzf99MEbkux+jEW+QsNaPhDitLWlUuiB1sScPG99PVX/f1vI4XmypH+G+6u79v
lMGg/gyTp7x0Np5yq/jqds141Pi/p6gOn1nH0Je5UpELNUVNIFaKZrwp3/7UTdvxh+/AMtegUf4P
gqHA4WyLhAov7S7itFnkY2IUGB5aFzYxYTHGABsFy+bmBmTNqT0pbaNSVsuxZP3xPtfpd3guNkE3
ChwaTIOTi3eZRfMfS1Ckclyz8+ojZ2Fkgw34nrI+iQDmxvPKKxyHNVdv2tsb1OpxrQ409K2suckf
WYPJWXvVzbjur6bamtjEsMa6gDmC69cPvEu/LHV6sG6MrdHl8/WNPGTTyoCxWFjKivnjZC98/Jsl
VRY8qEjFs+M359+J0cDzbtsMGmZr7pSkc5yWAWOH+b+1dkQae0+uPnzy62WNHbLYonmmnYeB1PXE
pcx8E9KSD/npnkNv0kslB3I+izTk/Odkc65nr5FVLmhhDTgANqGqDUuTxA0KL1pgiyUfxFenWsa2
D1/kG+qV62JTSfz+9fmcDbsKoilr8eaiSFN7+F2HVQLGJ3oBOW1tyh6nV2cCT2M6NR/JFjaZT9mm
IutdwgIm1XhayBW27vadKljzx8KEYyn7JtUxbqzg95nPXNZFEHxskDluuXzYJ0hokxnx0nig6/Dv
hN372zt///FgyNRML/LMWFioNqwX5W4mG2cIwfY4+bczafS107MwmEncNMozsTV9N0OfGoneNFFB
/ImOfKk61H7NBmUJc5mADo5OSMO1rRB/VOKf+v6IrebayLMhgIZkuSntEiXXNZ3KkdmuFMp/S07x
upK8YGvf9KXKagFmaHmlGBsmwNKXXP9kabEF3+mGreOyl7LSVk4WW9UsBRBiSQqOxfzv+h4JSDSA
IIbR40b7z/htarW2dJBctuCfC2O1TUR1ZSriFikCUisBFb/idvECGIImk3VPYZ3ZG3ZwAur9iPmn
bzCA4H6YYSOP4u1L2S86FDYk/dngebK34iCLJXT3Um6W0dvzG4mKHLMQ8TJTnXY3mFUf7Am6DqJT
wWDDpfDML8y4G3Ges3cloSJSI4FGccnF1r/xqxmy3kqbIxwiSCozCVp21Ep1Vsz2lq8NCRJH56+Q
oCDJhfmJl4kUXF4/aK1/EhDKsojgsplnLrADQEENVQazCOIt8wj+j27r2h1c9lF0mkZ/kJuZW300
qfo/2CI1f6VDWCCVdyND9NfPtASomVahsoNtXdzNhOrNgSaVlmD0uQkSRV6X9MrSbR6k3Tjq44fw
lpZ+awmpLQUMDhiljgjFIlX+H8Ct00tML+5I09Oib83d/gzst/lXF2ao2ODV9XC2SSedC3WCHNRt
UEf6KhMbgw4R3mPvvQRvbUwhtckx3OQ2rtRaeXhKozMvi6N9rtbFAiEfh9iYe6Jy45ypfvjjy+X7
K6LqQ/SPHgR9suzJ8AE7N6lxeqeCZGGvdEU7+c/vcL/7wewivqwZYS+EBbHAtqSpuzgNlkXB+zzA
O25MWUTcfLQUaUFBLDK9gRgpkfrgc0GN8VheArvZpeIrV1CcbVeCm350Ye+YVCOW+1AEUldgmwOD
sDN/5yQ8tRs+eDgTQQf9NUaf1bXxT5oWIUYScT+H70HhfIuYVxkwsxRDqmyIdnGJaQP3sJeFiPPQ
ZjYauR5rlS7Xx6MjGsj7BMANyHfzdfEbk+7CgtGPfX933ULKEzogALhmM3CVqumrvd5crEgbwGzz
JHH3cWriGsPcagLM3uSIuwdwopQorewOd2VjyrINk2jmVplAMvXASnUPVCmn1am5IikPCuf9d68Z
BTki3RS9fW0ygFwEi3825qrzoMNpZ3whhvHvh116VA1zI1/xBz7/mEshlJY0Tz4RYBukG5BeHgUA
XCdzGjwZ7uiYYj1jLdSrUrwBkCuJ5FqlbcCsbHJYevRAgvdsHJyC3vHo0S1F7zZUECbpA3eOhs5G
DkD7dV3UuUPT/dLZ/AXQir7jo33+zqIddrpsaKVLRg1vC2DQimHutLS6J053FCDUCpS70Pd48/oa
QPBOrhj+eEkl+ythceijvOqTD/1RrDCqn4QrtBuxKaKpTGQmzFK72IkQ5g2Kg/uL6cvnVwm8364g
HXMF9Tmhcsend9sMMZZpJnOX5lOMFlBNlLJbdao0T7gZwOsVYRslZgqpSVrPjH+ZBYgXdRjs1SZO
TjOpcE7HQWviUWpjN3Rd8+5TuVY2COTIRDBHDEo2oH7oe2tx82itxo8hOI8DXr5wQQNnZ9OR2PAx
0330GSQm4wqL86PR920qbrjBrhIWsQozsPcs7WitcqU6DoyE9XYASciN+iYqcGchQqQJpQgSikMf
Gzr69i1wk1c2crVgTjtjIocB3Nz0Q5ZiX4qVW1lE6Ka97Qy06NlpXxT5/l0UP9p8IJczSyJ46YS8
AL3+HxeTEk9qDkWH1BOGVHZv5UC2NUE1O3k/t9Wy/xQTfNNBF/s5WvPcDvMdc5mB5nR8LKfzIPm0
+KQXRuELCB90+218OUjtfcajmclY4ec8sQ5G4rm3s9slW2BTNDNPhrC8Kzl88avdccWsIceoYjrI
wIdpreNxELSUrVCgtly9mJqKmwmaDOFYoEVdFuxS73Y9SlXqQs4eTwrfbVZwBF1wZYuixPddgTAy
TrCu61Ema6/IgC1lY2bgaAsq0OEKiEvdwf/SBTqp7KWsmAhYT3gcTIvMgaEQ7wBU6ryKTTBTIQ3g
blnCd5Ptt2JbmfIhKGCwaZKAAPqXKj6F1P6224n+QrEKpUYi1xZ+2s4OmiQLamgfNQAvVHBg6Bmw
xvp6YBz9kzpwAU9XHjrzBnU0ny5NDart6PSDZMczRjJ7rkrl38TytUjGQguxWkiVMLnlocrkpuyN
aVEASPMVCPhyryIfF4ALnS/5hC1GtfFLqdM8YP348pVhocsUMAEOPidtp5OALf6PXQfKdlT+FGhc
uSuBDLLH97+gJHYiE6Il2Pb5TZoEY20IMuvCXK0ESrQBYRZoAk7FPiKJOwfJmjcXDkEx6VVNRgqo
LpB3/xjukrYz8MWILdT2tZ1Y0HnVW0RvyYmzJF5C6hzWKvigBFg5SGXjBJrmH/Ah46MR98XMP1OH
yphKIVgu2I9GrJj9EDUWSK7kqnNchYV7YtDxCgbw/yZqQVdpvI1X1RrcEgBbFMnjoNsCq47QoyBD
o1acFH4KBxAnp80iXeLmtnZaICt7PqpJoFIqGvrurniZsMvmq0o3oE+LQOolnPwpvXgziM+uM5fJ
AkDD2/u/28cwc8pzvB+YE/RhcZ3j6JyxoU54zVvpzC5vhsljaua7YKU4i4AmOQqPvUkbrhT2fI3D
nhM+FcF3a2Ez3qv1BaIWxRd5rdboXzzrx+MTnA4VjomtRGTjAlYiHFkQULbaP7dhEJdSTxgpnxcd
vC7b8TSKI0tnd/ZvOUbHU4oHxFzAkuUZrNUUoqp8AVHwoJtOMUqT0ZsYQ1eiNFSWmQsaLFSFmyZX
qoN2v4Vcf0+08JAkwUYaa70XgPpRFyzSoLbmWzU0CMRtD63QsNRUldVM6Ajp9xP9jE1SfQ0GB9s8
eQ2O6ebD9BuiUKHENKqqrBmBkeOaFc9JyzmsM08yAeMfJ8XBjtmH5BayC9BeV/NpIzqwdCf4KK2L
2vqfiUbHQm339VMd1d1BU1p6ed1O8WznpUq1AgU4TeSO56Avm4bx8jEOxP1pK/qHlBQ2t9jupj7n
JWaQDSj70dN6BrEI2oRGlECmAqVp+zCltchEfKNII64DSrfJSmqGZ5YgqBCKmldOzH+JAyX4NWND
vA/wgI1nx+2bd7vQemKWeCvlDzWFDpVaAOtVgRR/a5dGN3YUEBtHDUc/NRbQYuxv2WOSC7IZBTRW
RDdKU5jARNxGWNX9zMYPHVorDSSYgozp/1aOcnxCmjRWkNO30UZceZ0VO2CuUfy7yMhacLWwaNrI
g+HHcytuYdnL25j9vsTK4diqD5VrnJ62S6vwT8Tuktv5kOehjXGeX6Fm1zNOz0C9OKeHY0NuWUAl
OqJLY5jgmAF0hyfc3FH+hv9PJ/GDT2puOmXw5Gxu6rwKzlQBzgTznmhFQGynQn3jI9We0ykh+Jwe
ekABq6JO4/5PzKXcPrfDZF331w9x5fHYOwyEvzaioe5ZDiDW7AsY6fcvFQj71zjdD5503ScPzJpc
CM59P7fMRDUPNPAgv0AZ8yrEurfj9p37HkEsjaBop5LloecjZGZA+rSFCpZHqkajTyTT8qwRl6VJ
KkquyeVqP7+7afng6F2yHfD9RgpV74gaKOkRdwHnD5nZXMouaT00O68C2q9SkK6NWkMiwXwkWRKm
miR+cKSza+GKsozT073ksgHlorCj8z6MwTnno+OjaQLlUPizpoXI7VcUyTBMkEKQExxSRTL39aXJ
d6YxHSfTMjVewi9YYw7mrTE6i6eDp3xuS0sf33CsZuRJm66/QRhcKS9bXRF/StWgkzczREWgPUSY
ZYTDjzijoz2xs/vv/6moXWHh6WS0TPEOJCmzZy8QBHI1dQXlI9mRM2ruuQtGt1gTUKnuKFp+Zp9a
p7Xb9f+GTCjnVFhkqVzxkm0yvMn+7JH2OKrrl7Z9mJtrzHZbfvs7NZhQ4PDf/q6hnXXB/oVAjp95
/i/cWzP4SqF7fFb8k7t3iMD2RMQFjb8gi5Ce6qpMsiwHi5lFTcpbDNbVlJn/44G1POY+3fOWSGtX
NRUUMc0edn/EyXSojFWmKwxdXytg1Eve8OJ9ffmo2I831nzWbRdzUVYbVVtpJKNu6hdXEHm1+HSu
ZZCsvckwa+XAzCp5fSZfRGuSSl0Wq10iZnrlG0eBM5qBD8mxniqTzCsAul8oOC5NG/IWGktQ84HM
JaLwgYHca0TyxUd45ZeZdY8F96ixUltD9515wRvB2lYSqvJqsbgOcjR2NGi7lOnWQfoplkLBI3Qb
gGHccHLWQIhlZdeoCA0MOsMAysB5yba9NWDz6e/8Tf1Ep9ZjVU4PAiOUbUp7E2gLEaEQHXUI0QPn
CZH5qrKWLN9mvXRwZslGDNhpQUepV5PCz0xKSPvvqAt7+IA76nLAKf5r2r0YpK1JnpiaXhQovhnv
AI3anzIx6glTJdonjgV4aZEzqsepeec7Iqg50fWALClcWBlBoEJM0P/w7vYsCqOPY2VeI4Pm6NF8
YKJMUJrfZfGKab9CxeZirgsLOAlZAMsDBPOK+bJpUEfsXo56reGFE5GgkrdUvNy4230lDbDV4k4w
QpnZuSVJLv7VSZg137vJy0pxroB4cCLnRQHriy5ws7Zzyn3Mvadh1RwjlLLCU+rGlIbJcSeFRf2l
HleiUEY+RRKGB0IvnM54i5fMHqq+kCNCesUyZJqam95hEkFUSUt/XS3zZCc29jFCtyNpf7qO7AKN
isJvNBKoAMu1w3xqSvZUzmfk9j601wWRrERK+zeDCiTpdVpeYqgmbip/p5C0rHjmk2sEf1l92uNc
CDONummkGw5NPWa9zOkkueatEhLV5gotziyLwX0xe1m9WTq2NhXRQqEL1lVx9STbgRU4K/0OJDXM
EW1RhRnEoKakf2IDrMZ9XpM/8k7vOnrtGth0gct30j1CsdqAu7OTdfwPEYM0v9MeYxg6l8QOy7cq
+meezw1RhB93/DamZlt1sNpSzMTPyH8Bi4i7ySoAY12EIclw20wNzDJ4b3gbWtsuqk3CVNIZrHp4
XTbQHxsClofdSO8i9vBfUVuEQfKEb/FVWWMOd21CBQ7lZhVjt8CwvvECHcTlzm0m34tt8bRa5Wuc
jee7eSMX7Afx5XGnf+JNTpSX+AGKTs4sR8ysNH2CwHlLDeDBSEXT4ts75wgSDNAhoxI8CwtPSnr6
4K+qG8KH3hbXzhvj8tvgV8qs04FFlD9LFmGtwQh46N0jdtlCra8wZXgvmBtx4tzeKGQtxIxoO8aF
lggcpGl9kiaWzvBfXknnFKs8u3/Og2+l4kgwngc7hb4ByrMQpTa7Er+qF/Xo7LOGqFxQDmC+tjNC
1mnJDj1K6X5rqSmu6z1cZNR3lQS5Lz4xgjqEcW7exKxJenWGm7Wbh/NifRItMF7bEJG2nCeCzji/
vR+eJ+zk7MPrU+Uxy26G26WjW1Vbjfbg83oY1gEhPeM9AQI4IKJOcVXOIJLZ8dZ8+7ce1mVGxlWr
MdpAZL/DjFwjz1Hegcwks1+j51ScLbKGo6vDJGui/xI0d9FUCNDsXsDFJmfEesH+G+8QNZj7HmpG
eXWSv7r3LtEduVw8ZZNyzofdNTDfX0aCuJHlVtHALXtNnjHmJwniL7cVgv8af7PrZnDO2VE7dVtJ
PJRsn66zrI668tqwF1fbY05tMyJbFvlWPLC8i6fQe190WyZmHGK81H2A0diqjewK+lZsZNnGmjRM
Apxtz2+qTpQJUZbRWql0/IDCIUI5Z634wAVuZntPa4wDz5UiOjBa4FfxRVGxMZ7B+m9tYmGeGfkG
17LwQ5TAodroPwYkUpQh+fXejqR8U9G14IPVWTFLhhW4o80DHkNSm9B3RpSopTT14w74zIKUCs6Q
/2tbpbqSP0K87bhtHmAKBwJGBMgfIEjspzLbObU7bUDsaZtGF1/kqwQwtJ8hMisEtItVuNc0G/hK
Le4Z3yGNhX6fzqlLPYxKWVLlxrOODpPjaVBYjAMeNIn6UY7YyKc9Yye/5p6tpktAgvNRrkGfrtdn
/YN+ixxKNmZO2aLqlnZCZEFN0JeyEnvh/p/dtZZxgU61hJUJw6DZjluRV2w1UGnRiKOe8rMFxOrU
18TuKyhb+/GY96svPc5cSpH9bgtIoyrbrrjVCOYaaEDo+Z52PcnQ/4XE8fiuP/8dCU3boCnAp3by
lI/AfIiKYIpmh/ua9urkQfnxxBOGwBFkpVn2wTnNzJtM/+QQPlcNiAB8k+J6MLOQ69D+vNshcb+V
qiNqpr6IGFy617bEhqwosLvkGtCcMCl0jf3Ln9bHqz4qFn7dj5riTtqRWmSpZ1tjKzE+Nof9lIJS
nW3Q1bzRZXn7HOH9B7bMbnFSw8lQ35c1JBReYMIAxnxyei29+Xq8l6b4ulkbf54edxHHfa/lpaZa
o/U9YJNJRkJTqAEbhgpAkonpOdiShlEdubSZA8agBnReAOTDtxhskYCSAwsSGaVF0hwiZXXN0J+t
vrrbFqwsdUz1rLxlZZ7kgh+N21vFSd4zkJNPXodR1BgvRQlYfvTPrm3SQ5mqZHae/rge6T+Ci6r0
q776H+SgfGDvEVK7wtjfBIuC3LpKz7CSC0YLM5btvKow+oqWDZt4G9IK2qQAVomF7rS/EIHq3ZQK
TVPluI4NoSyrB5iWYu5KdHSVdjAtJ5pI0J84rqZ18avMIjAF+qeXZUohlzuaDhD1sy6ZJmfMs6i8
fZbEHJ5yeDg7UNhcbqt47WEA71lC+1AhRpSE1i9PwGBFS3Xl7TyafEydoXPAzE7Skx0zIw3xJal4
InqR9OITx+PTq2AZAMlS8W4eML3oXtrSxMcTnkgjQvY3GrqtgMg/8dVssgcnwLHd4eXABySWNUxV
0CFhR0089kfxXUIW7o6tYcczrywJ9qx7CxVzPMoZorW0thphCVc9LX3/hbbRIGGMkQatoX7zTdJC
MTxnho9an4b+N6/ED9tdTdKZo33n14Gyp80MVbderFZj6U6DjXfRyMo7G2SXHfKnzKYc8Zpzm7Vb
agcb+t4W7Ogan6oh6jxXNQpp3ZAiERNSxxtszGUC2f3mXqUG0WHQdkEOa1OpYKNCgZ1LpTJedYEw
3Mi8We2NFhpMcdN0o5p8MJv6JfF47YnzNJn1bcbZose1SVhh7vFCLvo3RSHlR3ZEoGAAdcXNvdMc
JGPxhaY7qU2YXEzsk8jxtVw/FFGF8U/TSUpFXd2Kjin2YQJfCZNnbgWBgduQbmXYoRMLD9zh04Fi
fTuVMStQxk2JgJ/GIqO0vLTBzIyTbvVP3ytR+ewxPPACRMn0L9d+RZYedBCXkhLOvj82OtgZeeFG
M8o7TB0o/QVGWQMaTH59G/LAlW3+CAm7tdWH0uCVGwc2yEfI1W17eGgOl0Bl6abLr5MZisTNPz+z
miNbDZ3C5fp3VqtvBmAwVfqTuOnTIo1ONrxUv5xx+3Bg6ymfnBM/ILyiGF7r7rb4k0gkDDZGKWpt
lQdMkMyvQqTig84wgdTRS/ldxAVyl3BLpDlIv0rtTfidSfyI0HFjs/GG9rtb4At6zqkAerFd6VnJ
QeyHAq85nINqD4mx2+jBkl4CQr8sXQtETIu3CpjAoKiTX4P8OJZHPgkvUPzX3yKA1ImI4RTIQsbk
SnpeQYiJB49eYnP7tl3zkpZbu4jAOHk3yxP0f98XTbWZgP2xckxxJr2IxjDQBOwCu9qcnpG11YjX
/6+q2h0dksA646YYoznzQUBVWt/UUiybZZPgPIWrMde8179sWCsFZgX6HDxxxmvf6sCsvXUJIXu6
gJcSzLTQTO4UbZ0ISChWhb9bHhazY5VKIIrr3bGkzKuQ+DX6mnO+RUxFAB10bEHpRehzUmQM5cIg
LwumNj+p0o/TbQEk8kIav0GG828DeNkTfv1mRVYOvvn7qh2RlyQJs6k8Wx/RuuqKDVbH0sngDy2L
kVZ4PeTbGb29bGxnxhs/WCG942s/zABxpALz8mA0w45NTBDmdH6lx/mLVMaRPRWuqS5EMykj4BP4
Z1CPDH0IZPOuJyfi1etc7FoGx5LO16+1Nr8F7nBum0MI38zp+BPKuRE+As8k8RvwYfkPSSxzqRr0
Qpt5hFbtQ0mKkc/IceObNZVWk7MHH4MSpNOQeh/6iV0fJl0Nr2fuvNCzn9eh+voyE5d98OA/b5a2
XZoGeyVRdu3bAifuJS6q7wKsZM9C2qsqS3KTM91JI7XHXTxoMmDMrmHuefs84Z/qonPJWcxhtB7Z
zpt92esN58yZvRPz8BMKLm+IZ7fSIE27H3XtHsJoV7iV4Lzosde6RCM1r369jVA7bQOUfCCQm9qA
dROe9n98dkuIKgClsusDVW5LL8Tku/51fOj5I/ewztH4EefuVH60vSfCQQfX/3KigmuN9J//M0Is
uohtoduONHerc9VYBGsCZkbCxBTOnPIJBDDHra1KTEM+6P5o9Zi2v5wv+G4k9HmEoc4yisxdsTkf
2+c3OD0t3gosFS/DUvGZ9E9ZNTasKSOtz8CtDqC2BZqEB46cBXjKdr/NgLzHgWwQ3cmu02jd/Rhc
i670ZGKSddaxuzeTW8wqc8QSEieoqtKnxcnlSw+MbRgtXZxPZ+R9MHsVkRFpkax3th6SO1+jjyBi
gwr/zPp0aNkMmLXNu0TwpmQmNGD2BxYh47Kri8VhzbL5EWzdZH97oxOTBs5rvVpHAUf8V8roCRDh
+hk5KJREehgYg8LXmpW+9TdHjtLFVbz2QqZPHGxKV35TcRwdYgplv2ZHVf1Cv5HT3EcpOv4EsYp1
UN2o+XZAoTPBPa0BTTmIHMj+/p+pBQn+h3mXIOZW19Gk8/gAU3DhJvLCYV2TEt8iyYqFYgX0t2Jp
C1Qsu64MrYiY84a7jFMD5+Xt5bXnvJ5DpaB1uCpX6Tc+9MSpca5sCiSvStG6TYaaNsYIuvRQjg4t
5Ptf/hRqwZDT2YFTYV0AopQU5O8bJZucDUgci0dAZa0fJYMRcZdnrLomlxbIafg6wUVfolfQcY7a
2h+oJu1EyEGR/i+i84nuMW49XWclwLThoH9mvuDEzZgwJL1wUYyWzwG02sNV8O7Yx/kmLWUII2NA
stitrRoo4pxt70NO7ZcCaLztSQ3QKr0nr0tv+HiGDdrvmT3jyu/40+BkDIvq5Abu/NEPWjH6d3Dx
SikK77byqBRKjrzYUzyrXeNJxH7d0ZYViryj5hfgA61eDj4vRnZk/DrsGrKanulPYqxRlzTWIrSg
fE/vaXjUXny1MduX2M0bgXW+2rgjAAVWa9CsdxwY1rNhh8lX6Obq9Btoo8F6tdgd2NBHPlWy02vz
3MYl8L1Mm94KrwhZd3HeaWGV1ijAOh+p92BOT5t3f0nEOhy5td8QfRXOtQH1nYgUkNd/JVHXv8Rn
aI8zR7J9TqoOrO8XZznuz9WSKr7RKuVRIGCPX2/WjqFN9KPuDeVgCUwmYWFq8cXNgZK4XnbbXkFD
DG8gPztqJTf5QWv4tM5rzBLvLPDKLQZ4FkvYhqGfeUhnYARnGCdkOg8pkNr/AtCk8GlEDeBsfW/u
UmAs5m+nI5PhwfkBKwbd2jaDaFaJ004jDuulzWqL0ejpHnYTssdabMWtq47YR689gQ23lY3JxXUi
UTg0bt1yuumMhFYW1M4XlSUXiB7NdKUIAVhrHEahAMLqNNXLpMnSlS6BC/tJ+BFoiqrV1jUfqPhg
lY1wkZs3vYr4laughHfesdpvuhtputJh8d6x4kViYhvL4aJDtYmb77j5zcH2jIBY8kxOZiI+kuvN
yBPQPADhGkYADA5iX0Qg9XYlv2nCS4fc5TvA+6ioAsM8wGaNAg2iYLyQoivGtQbNyABbUGOMCefz
LR4uhYurS0vTLOsz3eeJ+UmqdyjDjdsvW5Tm/WjmjFq1kDFhTQRdZgOn8BrUV4vsdjpLR9vbZ9nB
YCtwGjY348qUHR30NZ4TpzhoAZys7SK5ITYqm6J3ZT57ydcD3KWjU3l8zFn2WN/TnYUti0skE49h
iqsJdKEDIOnlG0BYO6WWcUIy+UZAQFkpSFmblqxvH3gGJkJ9BaJjohAa3G/daRU/0g0oVCgDf9dO
6Wrdq2NEjrKGvgpedHAruSFsmnNpLK2IPY4tYkWqnPlaeGvm6fwKrNGFpDPKmrQ8r58YCrisp/um
hGmea2UuRa6wMv10os8=
`protect end_protected
