`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MZ5EiNi8wWjejoOWJngTcI02I8XA/Tff4GDxh4Nhk1L35oJm3JqSrmAPvDE8+tFyYQFcDAFxH3bF
839DVeQrjg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rt21bsMFGBAdg9v3a3v1S8VpHfKIs8fDqMveUPyL2g/UyuaBLBRUvkEEhVvYJ/cTbB0sz7+Bd9cs
VZ2ceT880/nngsNKigdWft2YJ0a3tFoJ9bObAwuxOwjyPkx/q1V0c+0ayHNZK9eoOoQ2bzshHOBA
8p2aR22MsgbfOSoV1uw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BBIsm3yekMhTgZQtPuTz2oKTzJIZdlJ4Yb0GDFAZbIAzonZnDtBy7gPcQLfjUpByyV7isZ4H6khs
wjVOfmDQSsDjgileniKC3L+C+H5Z6dQ/cU+LHF/9/e0wGgodlzz13WLeT6vG16On3mfYKPDb78a5
C+KrkLHahxyp3PhgXHzZD2exrQSGPGCHZqL0r8FznOz/unlDEF11MsYJWc7h+FVoeyMApBJBnp++
JdUlIl6sf1ZDc2bYrMs3qNiSm7vQ+hC8YgrVqCm+rqPdMY2snx3M6bQB2Z8nGum7B6Z1D7XKqLa7
66rjqTHr+ERgVvAT3RBnkY05SV1Hk14loxeMVg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fzPidCQ0ZzS+xg2w9mSIrpgx4TPYgfvh5NcCVlQPjUQ8jXptS/ZAxY/HOAX3jfZ/evtNDTMdD0ds
erpArOFl+zaW8DzxOYRnIDDyDWEBYszPGc0xL7JVB3nZzhM3pC6+2NXBn35GwRKbqMjIIxcT0A7a
j+Walgpu/KvWwLkd2hE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IFVhajnFsHqteTODkUw6uQz+LM5uMDpwIGRo44Rol+OeYuFPUiPs9fOzBRaOL6EgG02H0s3RO+Hs
QKXXPbotiHvyrsuh6gp/+1FEiP1dKqDChOSc4R2CymTi65g1EYqKdRuUAAZmJ9tp/RApGrEOZ53l
7YmizZ3JHsX1/HJpxY3TMuCKwq08KMjcAjpfC9JdPx54XfHkEyGMtFphC9PVRKDwSMQnz6xZEkHZ
XFRD8hYNn/wKiPQzBPzzNfSLLes7P9NzJzS6PBijdaXYoR642B2ax181RLxlbTmllTcf3zetuSfv
ncWU+7wz6BxLpQDH6OP76hiAZK6Pm8pPbbW3eQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12592)
`protect data_block
4tfKwBzmD4hO9jQofXJZ5LKrwnUQ4ATIwxsjclNLPY9x6x1vTcp1pp8B3NtFFJGcGdyTjMJxL3gf
+OWxKEK/BNaD7zvoMsl1U5hriyFEtNOObHaosVjhu0zyWgaCyNQux2b78Zk8HlKIHiWey8d1B4j/
QXKyKqQPpE9LUpiKYDauN1BsFOUkhhgCdw7cmPBRDRn1JDyTACqkxLlzuIpvc1UsWAOaCQ7IQWpl
AyffJNxZ31Y8c1sR/1UBxHyWpPBcqPr19njjroS0h2oAwUbuVsEXY2P4ihgN4/zgpadKJIZheMh0
FZCCfKp+KYW73GhPg8kpOrs7vA/mlD8BUDm9SRdm0/A40IryVMUV45rkyZEUPxharwr/8N2ovW8C
1uXG8lVamzeG3yJAgv+b4NsXCcg9jpCo4utEXq/zsuKdIVogm+javg/RhmADPN6SdHGqIsJ4XxD6
ZqffgJj9TdZfIVghx+X5TQVNo4bsGKP8NXMkTz7RbNjVCLuxmuPW4HybR8Sn0dcmLMlSXWU4ERIu
ufCgcFYeRlNsbzux5gyUYdLArEdpGL+5vuuVRGb+98Qi+I1GZ/V5fPlh0EWGQsvcgIivm8sV6XJD
Ypsy4bnMXslhEoV9uEiJfRFyEhhVZZ5KHvn+1Bt1u7JCuYKwhUJpf0fu6HDuNp3HifurQxpwqpXf
HIOwGndbF4fAgCPUFw6FXrdAh0xrChm2ZNFqjYJBDm2L25lTY+vmgrYvjRiumrWmoeawS9bovBeA
ToqKvFXWX4qoGg5mnZFWX+ylv5u4QdQSjkPFp5Mrl4/TUVZPVGQ1d/6D5hdFd8X+y2EcY1QN2ehp
Dvx/PSjnbq7qyEjvGh7YpF63c0SR5oyVYbKKgaST08GNYEdj13uppA/ahsWuPHGBiIyceu0f2MAM
YsVgV7hAT/HikVhWBx8z5CAAi171AQ4W9QIVP50mOP0PMhrMRF6TiM+eJQbeuzwrAx+hN7S3a2FT
Wki7yZWJABBWjLKLcu29DEqjcQW1XuvSmBct26Y8emDmy61D4tix7Wdr0TKBtxRHTxmurlKbfRko
rLAZiCrpffv4noL1KVLX5eVvPc5UdOGfbveCHuAjG0sBCduGfFwiImkK+gVpAZW5a/hpf4bOChIC
nq7pfPaIVwZYkmG3YmPcvKHqEiGk69HHuMvcxSsfsBDCYg+pyR6yT28hjaXLgleL+bhOwjTTb/8b
oOENPUVeb6dwYPA7rcFn21peiAnhGmDW6tj02mMF0aaPvK4ThHjwXqiP61nnLzDIseEVdmKhJkVy
Pc6t/Th61nc/qWOZ7/CSCaJIrA/qwKVS264ZLss/mJQmrVrEiRlGTRgYxnqMv7oxO5G0ntjAmu9i
HH5ocGLvJcz9lCFy3cwG406thXNSU0DpHSDKhD29FXkI2+Hj6RpBizajQwhJ91wWvFT9TYJQ4zJo
Wwn29NCGQOKF9mMVLmZtGQdgUs45El9oSyLEkHrwPauEmH+N8g/sZuU733WSNL1B6/UEJdhQuFc1
e2+mtX1jPx3fZSnrCxEWXMLE6frhssjq1b8JAQXJ3yOk8sdJFlyf2U16qlEd9ybQIBiOr76UpeeC
a8TBq64SWzOVXRiGpBJzRLNpBkpxDAPRNZMXhZcQdoKg4njnXv9QqxfFkhlR9rT7KsPTrDnjDUaH
lt+bUlkmHAT5nxF3YmPGmal2C4Jn6YT6bB9appVTVLPAkRCrkHDYsXJgqEYkVqLKhwyswuTXvOxM
aSs3AIbrflxRpvnU/sLuskJVjla4CTSj6wuQXAcN8/SCvhu4YMaPJz+8DK15xoo7O4WFlyMJM9xv
D0j78o3YYMtNb8Aw7YFHm8wOKKz3mruoGkr2G5rvCREjw2A1bTHqYG3VuwW994A5/BK7jAByKa2f
9UUJPfXnMhYQyYrT9x4uDRt28jbruC8NdhTD7o52XR/skytC73q5S3XqH4evYKGjciMNm5q+BKfh
Kf2mvRs3QryS9ne/FQW8bH/ajsTQl3IMcujuCU7ycqblaCDlu/L9lR6sYapxNcos1dapT7ZAu+M7
Ssl9Vmy8Jy0UaEjrwz8xFaC+ezsiNjcdSt9xm1lGehfCP1F8mER7xzS6pUISbHEJ98bDyj2Tg3yK
1ZKbKs0aKrIiJc18mDlsTDcGLdf0dk/QLflB27T42HzLwUauVOgFy+EOZ75gaQ4F8N0nQU8q70Ti
NGIg16tXf2MRnRCk/ZIY1Tatq/NBT58mS2XOwqf75KxeA1mNAx6Z4djedc90JzczIIk75L1usvwi
CocR19RcnbYeOat2MYBvBInGlDVDN+AS+ZYlWdnsZRBnQ49zVNipkR8N1iTZT2MAw7U7GZRaHlku
6SEBFA79IyY17dJoXj81cyPpTEaQf5+bxgOWyqwfsOpr2mIhHCrV1mNFzJ61Onjpz0w6gurbEy0e
WCZqXEZgu8WBfagRyuJlu1mmuE7J9meyvxoiwQCtf4odrjnI6Gy2X4ihAEpjQNFPQdppEJ5c32A5
kkmWFIC4XPZDTNmB/poKbetu2YRSaPC4G0iGbLzsyfJ15CUWcs4pAWqkdRVqNFlJQvyqmCK5ZneW
z3J/u2QEBFzwLohRJ+eh2sMTlQ5El+ckNBNo6k4Jwj43dIeGyaQy1NaJktY5CblgtcOtb7bICCay
81xJ/uD+o6+dw63RG//mHlCEhh6eq2ETpd6f5C8+aYc3nbTKd+kVBRgD43B0kfFH5tbPvgLVGtPG
DYqdjktZVrReZeKDEndaiiVwzSc4irXevAV5FAdwJVB2Csb6kqlbqAitdgyULN6LVkg1dY2HCgX0
+B9wDBM0KLhLtLTj3/Uuh3VIrFUmxaPRiWFtnCSpl1VF7FHdOO6yVz336zwqNDLG1cMgBSpGQ0MV
fnksW8PPo6pDVMm1Tl24a+01fj5UB+czy/wN5UorITL4QgoNAPjV85JKUCx3F4EGxTJ8Ve5EsaAl
lugtvu6j1FOQ8lrLHheaXyaUB1odC9lVNaxI/4xxP1bRKikPNLAnXdC88bDEzFRD0w/39cEEHz4k
SwnX8DYA6R+m5dhvOGRNXJY/NgKqv6ThQJv3mhprH0Yqj0PXAZys3Q/9YiqNjroqKHGkgR7tDvfJ
EzIsGPX5myoYpLcs0l+tMnu/0k3nU+xyg2pS2JQFIFCIn3ekpaf/xp5PCDPr4vfKMRa1YWUjG+8o
+P2Ca1ne2MoyHhWBfCRINML+7pdI1eO+myWuqVv40oVrE+0MLIH+sG0x3Z66B9A/actHcLmELvwI
jiP2DiCwGgxDGdqZVCG6+m5MaCB20MGzYz8/7lUvC0I7lgf2Mg+vnkNmYDpUf/hIALvl5E1VhMIe
V3jowXErBsSZPQvBj4nSqPxdZFie4yPw2IvYs8fYHwBjEfQFS/4SjbA81bEymIuCGg3BI7MMY0yu
48D+zCFCTqJo7+iMytifh3rmbGlNcYN/i8Tx6tgh87VdPaFiQruCVRcQrPht7DLo7m7tCwU4XZf2
QKHWG14ul4JxFNuaOF5jAb6f8LBAI/EFG06VgQeuBmFSdCR2Oka79/6+K/+M2uNXcPIjdcLAX770
rWaQeFjW1VaFcKuXMhgP0HEfeULiWLXgabCNLudOgYqRW2Ll3jXOw95k429DsZsBL61CJ3/zWrlY
xo9A1epLRx+Ek7/8XgCn8/YkNsfaZrTn9qxuPM+aW4jSTGddHCt7AP84geeNWqI+2mkj2cCGSfIn
BpIp15Gl1z35B5SBHJGrT9SWKKEvXXUQ9C7T3mR50lRd/ifHo0REzXRbDXOmk55fjdjov+qFlz36
wgquhULhpca12mGZ6K29/621y4iAW5Jk+okjEgZLmT08UQxI84+Uwcjh6plNRuXgBho8oyYjHi6O
GkswO6RAY1YcJ+7ga/dtZIdaq92AtaoUOWS3xezuZ5k7OQMTu/ySqsteQxJVB6OJWQ7XRAa+VtiJ
qTvzDEwN1Fm0WIn+PaR/u8zOOoyoF86M97iaZZRYLFBcB024rUgdiZBs89r3qmdHcAYd0jOL6Zeb
DP8z0Br6GVXQBhIoMr/2U2VFDFqNSyBSr+5bUr3Ry1DqwWQrCRkJFpyWC/Kv8hYPUF0OBJ+dLQIU
2QT+CXUucEsyLtX1yMFdIeit6/oeKHjBIusSsIT+kfu3njJ9QfH4g4AYCdnM60meGM7xcZM66FXi
UcGlhdVGjOFO7lTbuQRUJHQA6XnajdG1cxzLi0W5zBx/siVy2RBP1x6QLG8kUGmRy02Zj0hlDRTQ
uM7TOiEYFdw6gDx5ZmbtmsPm7HO5nKYd1Q0kQrOJovKkJyCy+EGR/yTtpV2eOkUdFSm4AQimGOzX
hYIcopGZh/evTYzhTmM9YeV4AIy/iKSDt4aphgEpRkxKIeCqgdaCPPV7/qdrkBPMLh3B5mwbYPzO
pSBMc00YHPpFCs5EtC4MDsCIav++CawQGDl1CFJkTs9u1t+BmAO0QbzZpr9jtePos0rfYEwGqZKN
YHLVwAkLgetb+FCeBSjtck2mRFTsfeL9dUDm9X9SGFL8trdZuXugS2JBIujp9bMEQKy1O/JBj5Je
Av8Y9HXBuPgCm141OgRUZ0N93usOu6XzRnPs4r5bLGf4bfFm9JSkw4i31EL70njSEw5eiIuMgYVA
RmvZDk27MqZ/MdifHC/fDp4JlEwYpsx0deEVKn7eR6pLc5SJD6V+Wc8Ow8/PTBE4hCYZzuL9g7Vk
nOaP0MO/FZLJEGwuUEHNd2Y5h6AOKu0t1CXMFsIVV8x5Z785si+zRmwSx9mnIb/WVazztx6sDg0v
dzh8+QreIbuV4wx2G4UWDznIQMH3i7R89gymOnJ2H4LZe3VjNgM5H722PfmbkmN2Gc44lJK+Er2C
+gOcTmof5lRvENDAWGZ78e4JZPiiO1zRBweobWH84v5DkGvkKXpW14rntO/GX0LUQ2CfMbFDwhzg
iXbKCjb5aGEmlEDQn60mkPzMMq1PoJVK6isrcxFARZDdLIt/ricFcJGBVfv64SXzGPAQM1qoFZsX
i+DrpHydM0PG2whJNw37rFesL0+aRFMlPv2KkwlcV1eJyzFYtkqsG8mg09XNdCFxIs8+ctPQ95/4
+LmEmZ4L2GtaY2PStZLuiVW+03eA1QraNjcPqnzxGGs1L/Q+Sbq3YCmUJRWmKxHhulmvDaD2ANr6
0ZFOzvYP4lQRaQR2zs2+dtM5QOgGRREHjsxNp5isvqOvUXpDfoKB4nUUZJowtygmc/QEZIpg/4tR
4n687NRPoqNZqn/unHJ5uU59ElBDUfjkg1JvMDAu5GsbBzAxxDXB71Qg4vDgo6wlcAHjaD9EPFdB
br4bDvBiLarNVQTOYhAhHZo/1HjAL5N3nI9TMhg8XRnIF4LiEsZXZ/oQixuw/AJTqXJSu/Dj5Tym
Nz7oG9kEQikFJAewNg6euMp0WRXgzzVOWNg/RT6oN1Ep9tqWTeWe5tJIhlxghr6gDgHLQRo2HTSH
AJoewOlSlu6GEXRlOWG3SpMqJotvMfHbgTtIrUWpg8IWnUTWe/Z1XotUkm9Jsg/8fjvv62vYDG/L
nizNQwcFCjv6wqORzzAr3DCKFnrDQdKXXfsT+pH6f7qUAh4jr+DlaMUvEyTP1yFgF6yssB5dzIgU
kIXbFphQbkvs5NysqExG8og4nBvPNHviC3frUcsu0Y5upRYYBPUlWxbMKmGOjqG7hksiD1J3fTUv
oRmjbwuZ3r3XnphWQtIaxNn4fALCWL0NVwRfem55e4cSuA8D91a05lf6FUtHHnpjjNvLokpToQ63
0W+sl5WClmXFaLa06GfIDqkro2MYjdJES1xP3HgUTvVcx749sZa86+jg/RzBeQa16cPisKNEu3b1
jsJ/hFVGOo9SP5hF7KlCHPdbVAYl/CFPo7kSoH/P2AknjMbn/AhmdHjhWZKIHLvhpRaWXx9IMHcc
9JMRBdxEBKVMI49VvHG8r9pDBxS9tEBjYi7QhG4jefZVWkmHe529W5u167G/Un/YYieKrRF4sixK
VRkGCKIaMtS+sa1Pgce4rC2UkFoW0Yxx2K+Lejo3WIyJbGMIf32fE/zyqsHxtna2gHKORgZTpeIM
P3d+YlyKweI/QmGycMU/kr1KjqYg8p/VAk1x0J+Dx/iQp8SyDTN5wxWHa1s3iEWqrIKzkrLUj1IX
BPQcJL2jpfkG8sPyExmBfIoHTx0KcJSzGr5itb4dkUpwE+6rreVWGNsYcwygM0Jh3/PbQ4YIhd/9
A/hU724SSxzCDJwZu9JFwDvZqcKIKVBcf8elrp89stQmzhB7i+KuOJzz9W4DBgbZ94uIiaICQKwf
RPcmQo7QlVYnYP1u8oi20y1iA+qCwkL7u9fAwVlXgR2MadmIqAY/CtXYBS95hfEvjfrTIsiM0Nvh
tTSD/iQKS760uFBydti04RRuMRT1D95S7X9KTEoEmTxyPvuzgsAbJIKZjt0Da/5m7do7/u3ZsZ3U
ICJUf16QZosDC5xuBpZk2z2UkUZ92PWk0LFYGjlNZj0a0pzDsxC3KP7tcUrIQ6ZbBMuPDthg6H17
iV3FXToqV3apVMa/WWTSMlVEVZ6BntQpxcpCNg0OJ+WS3hBnLDN/d6CxyBLN2KFhPYc1aL84LmNS
G+ikijkEy2ke5zOKjPNsPMQNX3fKOgX8/RrhixJ0y7eSbe1FyqBt/AMCZBotkw+WmMkWijvUXXFn
xaRorqmXYRGpZlfo+a0tF012ORqTk1FTgfii7gmSOlXAgG4f8w34Cgfv8FkuFOSYQNahaNRX3xEm
KMu7aXiqE9PDXRNRq/bjjA6vEXyDIBTLz0zOGAXTLeZEGMrOaEx2PK60/M/0NPLYfsuWakxGXmHb
Rli7NsKoglbhlfdLPJCzXjlHpd1kU2xJbJHASpbpQ5xOrL5VDLXGJqlHrtiexRJwcQMnyP8VqfaL
uiq8lEg66H2Nbdqp4NHTUvW731nZlQjXJCaNJRTVQD889Q2mayOUcKzXpDabMyTtgwojKhZcVAVK
+RwjIPJV9DC5UOq8fd+xDbR5vocP9XRbBZ1mtIuKC12L0PXDYl+Pr2j0mjcPfAq4wYER3WBfMKkA
8qPSjVbS4xz2WUZ0zOuvDBjY+DYPgzqj/WcTdnmfHpIh7L2N+lB7Ah2EyViCkt8qXWjqFU65sHOu
r/OVSv1zf7Mi8Qo6YhKS1GZAWQpZrcL6xOSyQiD/rNwJGl8ApK1vKEeufTOl+iksLnxxgMIBNkiA
wYMUGaOGPHGEb64bDSR+phCSuTN4E3/Pg/PXI2KCYzEktT1//5c3F94QvQTW0YQy0lv9ZmxR1E+i
EqvPx/2bmFylIN0k05zUTsD0W7BOae6jiVBcDTXvw+2vsU7xq4DUYzbUXZeNUxZDzjIuBPE7afKt
xX3JFwmiZNrldsTwMd0LvfNvkaXeqGdF1l0a8x1kXws6BpI4tBy8t9BRkCsyza5ghb91/KiNOCvj
laXgYegA3MnZm7mf8OmJJAH5eS0pxDTNaa9ycHX1sqgLR7ir5I598v7Lut9qviDQf9jpD0MvsJGt
/bc1TaKI83LN/xVMN7pe6LovOcAqJ9uMQX3Cq/AI82OyC7QZgoYSzl4REnGwwnWsypSujFtnElfR
QRgKWMdP8xx9htJa3wkXLH3m3OYTVkRFlkLJCLxvZ9px2PiajdYqdELRmdH64c/iM3w2i4pCt3pK
OLmBCXLqZnvP43rwjqtsGwyIZ1GHalWRnllPcPNueDJEIFwwzDzt0/Ah6d74XCAgWbbcjcU42M8J
WKj+cYW414lJuHnfm8soGOe8vPs5bjHx0CLuhUnuknxsevWYDQvjW/Nk44pDrDldX/9VCJjjOn2S
aUFmpojrzpNqiSgmoQEbS1RnZLnFFvrZI97C9KAJxrc4AQDX43ykUv+soPGm5It+ru6h9x5+82nU
XUScD6C8/cJ4iMVaQXIEPWDpDzgsdYbEwleKpS1h1feg73mstINXcnMMtqDn1NOAXAvMrBefb1rM
Iqth/5uzhBPb7BfWnYR5l+EpkT4SrnadfNSfGEXFr1PFgXZfGd24Z00KNFa340LpkYMGIUrZo4k5
vCFi3+odgRoSGM2Cf9V6gpkI0/WD+3X7+vwlpB5iEWstyE7Senj15qxVXhD+2yq4/ka9jf8SiBRs
xowa1dVkEhZuTdRDIvXttUOlkRQS6DhKXjjw1dByhUGdXGKaJEGR7BlmMhYkrSWa1N2HV2DqYyDt
8y69004oLl3shqsrRcHFCmqpVIAu+PLkPOuEcz6oIftxnl9KNiH2kYGj0C4b/NnVyiLSU8U604jA
+ohHdhJIyoGMyHp6kHabJJvpV1Xp5J/qt+w+YhwC7CvHsz2VquuZ2uJOCsFlNwBA8GlvVXhacHlI
o4LYe7i6q1bN+i3dk6wsw4TSthknJIcO4+Ow8JQ+LHKAmsdwpz1Boxsv8LqC5HkiBGi8g+Y8L9i4
syRvRJoXi978F4CzWT35ZhrzaB/oq394wwKoFfIPFS92yqCGALJz1FDNWBeo4OVcwMEpAilSR6kL
P9IB1m7jceTrx/XUWmbcEetEpUEvganuOQYNA5sqhpd/3JKhrzwrBc5tMR67UjdJANqGjX4iGIzx
o80Wf9pHwXIx803XgPYKwt/xNki6ZmYQ/ZGc4h3FrBm2FP0U1EmMl3Z74sF8K0ceJBy9ejZJCcx2
kLu3h5ty3NXM/0P3teC/bki5R18FdBxXwv1iXTn+DbADddcWe/FjWllm1cZvAVCNW7Cr0fR6T0ma
EBUOzUynPoeg9qNr5yWTTHzd7iSrZja+79U02OwAwglLAOpkPe/ivDRw53oenvncdr27ReuSP6pQ
dHtN3xTVBxu/18ZgcUmfM0ei9+IclsunZ2IzyySLAHaIaLg3jEKGfHcWV5y7EThaXG9I7ETECBRp
Bb2X4x1czv+oWEeL9ZpxdN2D/QjMe8cmUmM8lcqdB7ZaYgWBHoXxvm7Wq2Ifk7cihh2EuiojzZS0
T42cawumZHT9XnEagAYPtV+URhrwYf7jcXUgw38xAgsLdRunuuRH1nbEbetihEahteIQ4ubo93GS
n95XAMgNtNR9BoneE6zmHJjE0xqXOV26JC7p/csyfU6ON/+LGOu6dmExLwCMBH/dAVRu/TpGKHjd
SQSy9BpJjaOB/CaXaZevtspa8K1kQVwOnYcSv1+HaU9rlsN+T75dZw/Q1qpMzN6jswopCdEmnxbp
SCxYTDSAWeNUtfN/+8vYbfJO96v9J+GtrFCmH/duSJ3PtOoQYQ5trbXAMLWC4EXhg9VrkvbCwBXJ
fOxGD9j8mkVEksyJfXhY5TbkoxEn4ZCGBkOgGN2tLneaKblnEf1YeFIHsrPSOlMSiyvXuagpu9gy
Yp5YVYUi5XdrTU+LXBZbIIiUWnZb0blEyRKSvAgnsQMFGwGbi+sukbVbZJv243W7Nw3EQmNxUYV+
gsJqL3Ubg4XD/O2WmgtR9RNF8wjfkoOpF0/XAKpOoSllyJiyUrS7gabbERipz56mNiWhRGGYVPjm
P14/rs/x0SdJEqtgzCkjNPk29xfpSqK3GXg3m1OkQdxlD/uFofXlvKzrXJDODn+E/Z+mknID91bE
WhzEdr9WlsTBeqgzZcfASpenO6sVa4ssUP53i1hiDmEx5kDrvODmz4uGPBVdTSg4SPzSU9kkDE0f
Unbiv0pBlKS3t7ciWQ+cbWM6iajmjyI+d+ux2i45KQcIi0VBghezT9Uhmgx3LldqvAFMcfMdtNRI
TMLSLgTe4OL2RqUvsvEQ7uvYPjPyJRTI4ErYFGo9pOxKVbIICOnuhqzl9P3QZL3Efu84MWne43S3
pfnKZEEevLdmQnL42685F2575HXsjSdWMQBpcBhHEjE9e612AtyHPrKeszOrP3ZYu5YgYfmQX/5u
w28x7O8voQnDKsa9IgZEF3UckozsiVaUhifD8HcfupaYsQhLE2CpCuwDnfEz0KOyR9tWXqvfysW6
OXP2UH529db53hknbAVBYJ6BRd1mM0jenVAiU0vOmgbNsmV1kZCB9dIOpsFBwM0q7ulml/9wqigl
To6WMe7tNijA8uFaFWHR2gne/kLkphMkfopSD17BNyS40+OfFDrgi1IY3UxCo2lyTjtnAQipC1DZ
QAVzMFoWSGTsmaWM5HeNBbJvt8B74oTcxpx7yyP+5bktPy7oSpU/GMdY/zcAOW9Sy5FpnWduhrDP
PT5qz/JcO3QGlYZiCDBhc2lOivqjUyQTffEuVB+euDyYJIeS0+gPzF6Lz4Q+iWoIHE54IH+68Qlb
h59i7Wrj+1eI2tjuqCo87WthsNHluJWdCODXcU0Nn9WjKkaXE6+kHHajKzOAUFrnO60QfpPvPcuD
Zi+aass1f4MSXRYge/s0Z58b6dwzwJ3wkuGF/rGJ1q/evWYPu/KxOvjTywesGuqoHaUsUNiZ6Yvv
cqyOwVhA3hvgn4FfUE0J8Q5s6+0Pm0x//mZoDpFscx7+/btZAFbp4BeIuXtk/XoVtWydUISKCK2D
a7u5LcloS1lCLDcss2QBFgHYPAsvq3K3hFy0ZG0h1rcgo3Q2V3BeA0o36r4OLzLirN3rEi4GPKix
KoTz80lJgXdNAQee415ca+84WuBwRV1ouuxswCm+zKSNttIaCQU4fvjUBm1/C350NQOVGGxJR1qG
+Dbi9+UXyNZ8MW48uw86ceBNn4Rr38NFbaNIpYjEmEhDc1oMeC1kvZoEWvBDu74B1zRiXD5UcaBC
4ea074jmiY9jUo8TTgnbP4CemQlr4LaItc3nAc4G76NrDoQAS2GTUixiAlMQc0MmPxn/FYQTB2Qe
AnwdbjXMtPHLPJKK4FRd5EOh11fXfaRTygvy0GcOSMZR7z8zkGEcpzVQitNpKHY1hIl5ogy51a4B
H9s+XfY+6DsYrRYiNrLWb9kScubyOBdXJDrFmlo3C4HhqUJlpUSOfPISgP0fKU8Vgln4M5zqR0Wz
HOs1wcLTb88calWl2XXzyTAGChVMfUqBkrQOB4LCRvuseKcJyttnvNH6lTY/PsXP2eZcQBJwmqwP
TkZGGn2JRc/cbhQHP45dOFbfWN15/uP0R0VTL8drn0OF6n5n3v6hVwrgpF9BDFqq7/HY0s55WRRF
glAfxTev0KStXf+aurCb85W7aVtmotNY4EqtH65/cE7FyPGGwKnpvDLBsFT+zNUN9gwy7pc0CYhh
/lBSXL1us4twsZtZo+my2HaQK3RxJNZl/cvp8LSUH/nq368b9e0+bikdKjU5xzG3fiPnkiXQH7tJ
/cpkFOzbAyE78PnsWIfPPRBgPYmAOIWya8/QX3y4IGwrxO0aBAexLakP47/0ukjbIxBlPa9iFRD9
EjYFpcTf6FA0UlBcKliXFsGDY08uRhprdmkr0TaTA/5fequwTL7M1golBd+ME6pSFoGk/VUuYICn
bn7aZpVt3G7N6s2t5bzDiU0FiOeWcjPbo94gKGxwGeJO220Bgz0gTQfGVigUwcfrtm2TnCJ6w0Sp
Q+zKy4VFqJoRrVYHaCOQPJRro1MS1/jTeN4uwjKxuNkiG4G9Dud74VIGEoCHXPBRgqv3R2idolpQ
REr4ljGY8jHCNYC/Zt+rCMoHkghioA1Gl9370nMN6oB5opTbUcFIlmgx0qb6oYHxYWq0hm5KV4An
Ac2UjFYBlEEgb0BMXaV1173bunMLC8JRucAgjiddmKFi4b7RU9lPWhTDPt5o8xZwDaK/iwoIrrbu
Kjriy7Rh/yZ43KDYtAMmN2Slth4W3NLXQH9oOIafVuNFVGXu/KlzcZrgDffUaQeUl5IMP0baOcFd
AjQJpmFuTJKbrdCWc/YXwv5lo8RidPfx4o99A0wZfW1ABaxruw5C1dAY/GxtBkXa2E/AH1zrD+Qi
D6AkTdhjGTDr5AVGHiN6p81fxkO1VLm5XCt3iozsYs2WmFzfKy5mTtOIWX1J+gcFta0W6Cpn4vVu
78PLHEcxKooR8SONSXiF/IGyLHWOXn+2AGNTnQcuBTRwqTQoxyMPzXX6lOqpWu0SLjgZ6sLs6RO6
emPKdtUlXFSuuwAT5LSJF9ZP26J9Y/+PhPJbBZq7x/5cL656xLZupXrUv8iIS1kRHATS1c/pjlpK
w38dRZMsdJU3hSVQ0cU6h8LaNK9em6dyAzRu9W8NT75d6UhtcHqdLVKEvVVuGwdilv5Xnk0CFKpp
Lcitb9obigPxJvMPHdn9N61I40CF9JrsYOpGprDB9L1zM52Wi0xsreiV1uOS63amLaYb1jS6eQfn
G6IqBcNrUSolGmNqsMZxgwnffSXDdphAcAF5MPXyaDZ/7vXKzrFiY6Wyp56H0BWMQDjL5wPvzvY7
PLzy5kKXJgzVUwY6WhO1t+bN2yWRMR+gl2DigDhd5ys/r9mnwfrHxJ4mYijQsTT6CS/ny736TxDl
vkoiuikog+icxF37FeedclOsrLIcBQgo3VzJT5po8lkLwGuCMJsTlAm9jmQFUxVrF7r3gkjkvMTw
JXLc2DtiM60Qpr6A0FWY7v3h3PFJJH5cfFLBomrms68w+piGQxZmCn9laZpwrFv9LSrb0MrKbcGJ
kf8ukWAJ5tv7ghk9ZLLVWCbbWZ9aekZLB951arKIhTqexG5EcGLBWwlSI6f55paXGHohs3rTua1f
xXMQswUdxJYMl6gJSUMOtxSrmIRR2lymIoe0/0r0QZIKxAemXBIPpA0W9i5ZSgjuLPMmqLYnuxFm
SThxjZT9bq8g2pa3RGm2WBKg8z3T4o4dEKr+FBCwIcZz5opzHPoHO5jDoCOI5ZW34KJaDKNLADue
3HuDic12MUWjXgcsCF4tOYZv9LnB0bIAUh4Jdql3sOzz5jD45x8YKfTqiUSqvVMAPpFYmyamxjjl
4o34TfbKHbC7ABU7l9o4GW8pdEtw5dlE2HpaokIJ0v/iOyiQ1WKdB0hjSOApgsa8trTdiAHOKh4k
KSslMU5vDOAO2LBg5o5ndR4Edk9O02VE2CYkPCLX9IWfetioR9DYSS4YUgsycNZUDu6J1cATZZxl
8302W199MzKd+6rvTARkyFo1cr2UIn8M1npce15TCdyF/ogzaFYMHx9pCozSNlx2epC9ZDR7LEUN
eKfBEDVudAiOLck1tn0KoO77oEmmoCOxuhjqjqihqR+P+A0YRdejs/uyGwZr221jVC3fGVIquCAZ
O7uaufcXE+iwpnthgDNBb8jUDb+Hk3bS7U+u3DjHE8SQX5m/OxNb/ZBhB/gbxEFW5wKQFmW9kdPk
0C6J/54ihIEfguP9D9Ivu0mispDQttTmy6OegWfc2g+9dM/kXaFoWGHbxgVrRZzzxFMgOTcqVoc5
QcHkJ3j+5caE72EFgAODEDLvNm7L0vBnrXKXSjPHdtx4TXLA/X/aiHrcex2e2KMsDYc/W0YRdG3d
KiH9RcS6tR3QoXGz+I2dUL+LzSzkmoFffcLQ9/YaS3TSI86iU5yMmRHF2SSWM1yvEEzM4Yth6nPm
7zgvkWYiKRHEFbf20wklRQJk2G8+X4stJv0j/l7Qqu3mPAwveJD1t79lOD+5P1jS/S/EiC9Lvo0J
Ll+70senD6RaJr6biJFO04LO57H0otoAg1G3CXJmEn/32wIhj5W0YJp1a6Y+Mtegh0ywJ06qkEu1
eQj07hwxomvwf9jku3ctQwYanaf9ubbjPcTsZp9RsMIDfYSu7W4U1XDG1pewi3sLqGOMpcC+5L0R
AT5vf053xQxqEphauU8TXAwUlY2sRbeChwy2GXoObq/7Dv/C+LjXn4oZusASRTHqVLah3d7NIer6
6xUQLAU/6thtap8+ofrEDxMciCea5ZoTr0Xo/+wv0OXFm1j7BITqR75m4SgXV2+c+4cN60GylSvq
V1Ci8FwxPmceJDfDsxRffwedzfkSksnzSQQeI2oa6SdwTG+LDuizZlSrYvCrUnJZbS/PZj9nAkwM
Qx7P8XvRvirPjBPUCVNGPdOncGDPv45sezCGHBGO1yn1y0IXp5vA2YE5MdhXe6WQNv3/CIN/4Vdk
n6swjYSdvb7ZAL538sSbxNIeYZgQu8L7bwILAdoNX1V4kMAHWAhKQtk1pSWwANLgm+7nCVm4nocp
k1cdqMyeid+WXpIZjldEhZHnvS1anYTNqVsGjAWH9XSBlVRmPBCJZi5ethc2NsGIXyISILev/yWy
lr2tAVhAkqeEoRofrVpr8C2PZzTN9Ks5vXqxdDB0z0SfAw+Ah1CT3ZnT6zk4bDasPqr5oRIF48Ff
mE+fdUKtdTQUZoo7iUdJu8UBKio3rQgvHq6t7FH2B3nrQVZvw9/H5Izx/feydYISlmvvEQLaKpjB
B+ihauvL0JrrOq/EOo6g/BVJhNpkqaGnlA4HSyPM7BrBXcOWxTkve0WXcuMTwqX35r7d6xY/TaZ0
MzgmWsE26Eh175O207bYGmeSIXXy/r8NPceAKMSpkB/XBV1X3VG7WM2A4nY3ApD5KryOwPM96a3V
RXxNs8DnkAYUO6zqx68MUv/W0pRqZxgncHESEetBXrJxEd1p7YjjIaTbymfBFog+acl/sRd+6muX
4iHcVjVzKKQU0be77wpAvFvP7O7x7MMddzN2+STTWHFPDOuyfXBUDAs6qyRpsaCRka1oVGT2kfuY
UlGYNwRCNfQ7qwFBHL3ItbBj6SWDN4FI1pmiqK+BiQu9sLco9U42/nCL8dlcpYYkQM+IOJPF0zZC
mUSh4VKWLqz7Z0/CPDgKMMZklIVQxtVyY/85QMq9e2rgW+5YFUPmO7ZQNfKoJ6kJ1F6uZdxyBvvr
GdMog5e5DumIuq3KcwCO1K8PWWcO5CGVm32briq6BcXzrocCHMrpWLdGXm3S9BNp0iB4SvBVIKz1
iU+2uhnSlfGokSYWE+HXFx1x3nrUwEfiXcw+xW51NIZFItesiKc8bjiZ6qHmsVx3C0vzdIC565sN
jvEI/dIMVhrpbuwBLn7o0c8yLcR01xr2rOd8vYphnrMnZ35IvamYLPzEJ+swC9P6qa1iyFRrjtuP
ULXQk9tQY3v/13+5JEVD/ykV8cE4Ouw6c3UwKGKElLLv9fgoPXEGEU1iSElJ8+KDat38NZcYPOW3
ZMIWkU1wn0vkDrV6AuCdOa/GxycjLewNksa508vQWBieOStjI7ibphY3qUPqoG/8/aj5R3RbcCr0
V9P1B8iIhUn2CkwAJFEe4tdOORs4roKx/NoN+wt+wz7Z+rZTLRlPfOcFzp3uS6Fefsw//nsVyUTJ
3Z0c9T9tqtcPW9ENb+sVGLfiOrr7XjB468mto0C6HaKm2AF5zlPgU5dCRWDfXKELaFlxolBWNs2H
RilJZtcctP9dT+6kSS3HvhGflSV7yYRB3orjSzumnKCVIH4e2rfGGoa/ZwpEMfkhK9ShxeXUeVkC
d3b73N0Bh+oZS1hk0AFgKcs6ya8vhmKKu+ihegrhU1/DXrfqP5TpZ41KwQjQPr5zeRZfsXmgIpwB
92SGZ7hcs/CKIs7qz2k2tozqOGxFk5mnu80RhEuBQ7dQgm7Fj5Ns7Sl6PYXUJ1a5xnNuBpUkNniG
YYQDw/7M77L9WN6kpqGThILhyCQRRJIK8dmGUvrkJw3QradQ1aoSLDWKccxeXJVT7S0BTgip6qQL
LQNP5DLUEoZ415XjbxraWavunyIZ7n+1NN5bypeCMhVHwIGeNaLFQDYv2t/FGt4Pl4sG5RP1k2JA
dfcUyZxWMVGepc4omc23gzrF2wCALjDCjD4+9zsaSYWoCA1t3i+hENfJcvvX19vk+7JZTQ4AsjJH
d2sRtFOJ8NNTc3CkeZoscVnBud/eC6XYzCklzqL49wUeqb9YloYPT2ZaFblnHRszC4EdUfctz/iS
ycw1SIxW5lMkIaOHnwrZk9zn5LoPRIx8X6FwYd4HgmV2lRnJnNGdgroERPcJB5GI/yOPPLLtg6ra
toFFkbyEX1PTP5uU58brNVAR3bfZPEJ/k8/RvBTkqtsTIJ31WbGGYgxVKSMnZpAya+ZhSZHvgJW9
FREkXUpVgXV7qhfAQtSoBsuEpBhGVeUehJu+e4+Ww6+iyL71T1Fi66ntxlhnE+92y5VkRNZo0275
s2EriBrvMxRqNKvps/fKdJIAg6YPZxOx+dD33OWmFgz+ZDZDlG6umgfr4U5vD4UctYluId9bd86M
tz9aM7iQ0sFX5cOUVBOzhvCe1+bimLmcbXxvpUB94TvmfXbtnstSovjaDyB3euNtaNQuZ3t8waCb
buXqv+BlE4FuhYbFGucxwyKgGBb49oW+OdsU07PeRzYpIxy+SwdjffC+n+Uk664v/0672NYPSWg6
s3k9j17avsYMQ/vUCXUgWcDnbIB3JFFGcmf04WTviysG9drlXzVOxWqB2yz5Xv5DXTfY/Vu5aJYT
vO12i0ufphjGlAKTuSAusYvLaPvzc0UWIwzv1I6U6gsDGzOkbhp3xIW5pOnWSOyDhzkIxIF6Dy+Q
9CzYzkJr238vc2jw9ADlYOtC+gcdmTppRC9UNtsnwfAv/pC2xovFjH/iP7MIricUuE8DCLciCXCA
ZUvrNkxYPyw+Cb0dgVYnBBaKAfC5Cu+B9vTlrz6fT2ddiUyW1wPhAug1yaoWb0/vlQfVgEStStlH
V7E3lP6/+QlUzUUGr/HmMqHjnVcq43+6cv1GYyESxcbAbJv3mepqMpUgrFWbS+XTyYMJHjlNLgsA
50rNKePak/8Jexm6TfMbvvyydzfsm+6DPmW0GFYfr282/2RLMgCHymN+get4Y3nItQ6200L23jIa
yZZ1pMhRGwFmxu+qHU26wSK/b0ze1CTwTj6yP2MuMGDMMFLKRRQLAPtvSTA2NrWGFMExGw==
`protect end_protected
