`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WFLjaaLJQKked8brra52FMrnU5gOzpUbYjBZyXcU54x75LOIpYuTJw4PVbEzx7yIdlRz6tSkNlNy
NoqMCrYt1Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GBOljTxmJ2YFZ0Ztk9wlIgq75eBl4lYt6Zb0NKUiMh3Gr5XBmfOIdnOqoMrc1GJ50QDi6XAbkNOs
5mn7wxZx95ouMWQJMHpZ2+yeE32ra7b9bqgKYPDaErZKqO5keH4aE6ljjcMumZ+wIZuw5uNekBy5
4eiOauN81L43Q1Zaoyo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z97wlqR3fq/jOtjYD4zyLdQWqTOghK2np+UabMDdBb5H18UB/MYbCf8dOrTvDHaJRCf78cI/1h6e
CXElnN2SHOWemkKopF++Wm2OJY+DxmELAH0EWoGS5czDJK7688bURdBiaD5QHWYgvKqrnPCvAC2f
0nyqEQLSfQMQ2tN2rbCLG4qFeRcDm6KqlaKS7sxSopNw51x9aT55MXIvhfNIpDjL5hnkrL6f+KSB
ojdsg/o+T+I2y95F0X07idw8XIax/Y7ri1bhsdHimPQgYryxux5eyq3BsKHCmDI7C+bM4KSYePyN
vg5p5tB6x2UJd+swyEkQD+GYuEXojYDQirhixA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aVrQ8ocezesdDOa3tVwp8PqVYDaRqxc+W7Dz/8sXwxd+MhWD7YQe1EliVcS/iUYKVctfQbNpCv0d
lpef4Ya7BnudWhaxGZT+dYVRgYvByssPmWJbL5kqqZtcI6RfjWHS/0wVGGpASv0A903YfbvaG4Ac
vmTzaapguJHHceKuJHI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ARIRhhKF68WRz4lMllQNXmUGdrVO2ZkZsTilngD2jALJnFbofjdqBe0paSYkQoARvDneaGcGvLcz
vnyM+ywA9UO2nKyM2mxrlU4O7CyFuF1gGRwOS0ah/l3V7vscGvY7P2dkTdpcxa6o0+MPTY9/xPX8
+j2SbrxYsvwrHU450T5UQfg4wlqDSziPZXttKXSN4sz9EuUVX0QGPmbLYysLNfIFmC6fmlbaPc+B
dRB78RaB4DMV0/x2po4NcLtRLur1Mn6FQ4w+9cCgo0rusHgIqLtpzneJoExzAlnhQX2NjVoFUjqd
/Gy22jcVUH/eFdUtzTiImGx31U/7GtW8hzdq1w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11616)
`protect data_block
zg7pO4GirxUiwUVLJQ7YYL3sZNjdtEqyQeh1yesHT0//HsbGYVd/rtNYOltxI7TQEM7PoluUFLuI
Xe8WOLeo1u+YEdETW9Qr9g88Q5sVpfPSrnn4Q4VL8CTOVeBpaygzebEvExub0HZkAZGIanyal3kc
QcgJYs32D1r3UST1thD5rIOZ6RYd9P3LRKvNjCyBOzV0DClsc+6I95ikNT6fqLA7DPHeetyucy+p
mIV9PA99dGyrYG4u2foIYHnJtAld44lJ1KEfZboFsJ1XSeSTA3vzTjw6I863Ea7hw2ekob1QXN+W
bjLvRC9Ma24B1IxKKEjpKDTUUKGMDw8JGNQpZtAOZrfNJLG3U6QRsPc++tnfxq6PCr2NE+zFuWDS
YM48ACTsfzu1ZQtd/dZQZwZqMPBLXg4xW16oQ0Y1qJjA7NvLdlyxgTlW4bK1OlKIih16CXuX+pUn
u/3bRXiPZMb7xtQvibRJt9xp/Zu+cZudSWBI1M2OVAYzw3Jmmdx8gQ/kmniHtmrJdC9eCsDNjDO2
K0sYmKlGXlQVqHAtA3k4tU5TC1J6uYAb/CJjaaAiU9DOEzvjGsIBbkdcgg9xDszCeVy4+t4MRLje
+xtfn8bDmywdjh20vlri806h44TMtNLBeoTFk6q5Z9wsHs8+5iU1xui60CFV+UBZTgcIUXjetltv
bzOAMr1WFODoFzP7OWzNrHq/pcNmHsIiIe30Ez7jkVTN1OhfviVwcQyUg1CNEFm5w5eNCL+I4O0H
ap+tE+HitROs49HNdAvzfs6Z0pzDOXyNaK4JrttGC3fINxPUtB3HOyNo/0UFufbCV8Bx2BnloULJ
F5/3jrGkwz5ClgYOJWwrhEpGtQ7TAKrQlry/JgEihEvNhjjJqInQp9z3lcceLR9s8ixLCmRiUGln
acCIOxfIiqtbnD+kxptXWNOzI9K5Y0toUObrPwD87ScDoo0JQXkfy3y9AwNIXO2/C21p0UXIIOHJ
yg1qrooxWJLJLEjs/DSiPPvB5CNqm15uDy7ZI9yNKfXNBn0H4VNsCpZhMxPEvAH/rlfOpNG0BKQr
DAsUw8PkKC+m31BrP4CDYj3KTMbczLJ81OE3Jtg7lzMMhwnJbzn1Mz0e3vMrJedwFrtdKcRoyS5n
01y07hKE6ZPSDFZwHLj05+a2ALdOfE6MmBc4hn9urdI6jDBv+tXz8VBk4okevfsImYI/uQUPHKkc
tsPdCGWdmT85XZnJCEX08f43GqOyluHUdY/u+fYLiMVrUEq3vsdTIzVsaGa6fPlvXdclFKXJTBUl
sxikWiHzv32xDGQJThVReXUTsMlMiIO06Xsii6rI5h2pVB9EqKgMKLA5oE5KC44RMU4eB8H92DrH
f+UBgAEztPJAdjEGduSDmtjwVlh2dUhNBSafFHjhbZWLYsAX+pWfAiHnHL3JeYpvhxbSyTTEPtp1
nPIXufJuUNnt9hcrqPsEA3xxq4ppZ2+Qke4xtDOzKi29s/Yd5swsy1pp/Iw7yDO8VrhJQIkVDNUI
elx7/h1S8jJh7/WwSpgZ1vyXuZPQdZ6aYs1Tdsjym6uhY2CKDYWf9H79xqvlbDC1PTgGzudoLMbo
syMV8RbWdySMHX6yORS2J8fSA8vYzlVgoMAstQB0+I01GxwdmxV+OJoXdlbbsGonDvpt51dXhtIF
oVoUrKg2G4aCgOA12l5rUmo/VVE0miwLRRSxoMVXDVsmc5qP9RDbqO1GydFwqn/WGJADYNgd3l2q
8xo3rwFmwXBStvEmxInAubu3c+JWLaTUtB6I9pL32MvztU/iUbZth7ECXW9ya3gsHlqUpPcGtQ65
m5xjLfC7x3IlSB6GpoWfL3iUvSYUDeGrLpNwFOLwFEtfR3PXC/Wivhd4Lr3bEJTxSW+pveJuR+41
x3r9J31ek+7q2ewoIxbph1YqmBnSWSndPryhry7Hu2SySjfh/J+SFTSkRoI3z41Xw3dfizMQ7NJd
iltP4clCOEIEsm8rQ+SbPp+nJk2RULkGXVorTgfAW98GhHmHOdtZZcGnpH3NvfEnKsIhO2e65UA0
vbgVb6Hh0+m/Vh+wOFaOHN4bbYuuAliwG9SBFjh3ozo2m7zhZ9uvyEPbJ45tEiJDZ65e4tyI5Kkm
WnCcGT3LncFz0SSbRAPVCjczaezSEPyCvRtEq8+jFRmg6Yt5KC5+i8IAFFsAcd/YQTb8mJ7Y7HEp
7QgFC85hz9tpGnNDW1EbGSSyNYWUshke6Prw7ZaxE6nyPI2oQRHtQkFVwchfiKYbyuomFdtNz3bK
pXSteB7VmPZJ7aQe4XMF1ao8/FM8QAgK1u7NqlxhkZ8mNVb1UkYDeWy/XOzcUodEyMALI1uBkv3d
K9IYisY2Ids6S1jwsooftV0iSVe3yfaFUWkipbrI8sb5Vy2+XlluRqRazY8/26KAcABx0Yh5j7oM
IzJ59Z7OACmdi4vA/3Oqxf0DTmnxj6oXelY0s1B2f8UXBVoON/u7Ppx/jBlnauifM/y7TDRun8hn
PpMJxG88bxhj7aLHKjw2mJ5L3BI3bG0bO3klnVJH5+IyUw0bYS1jHsF8rV0t0fOhc5GbT4dkcF7o
AyNzy6ax43emqC4D3HjSGHYyqyQuUT37hMrGKrHl+0I1n+n2z6ezbaEZGJetyUpgMC7hPEsX3Wjx
IOPx7870oXwWv9mhSIG3m8Xldx/4ZDCRO9tzpAUj31JhGILsVBE6rF/ueU0oQcBn1ncwPpwuIuhY
8BrsppuC3OOiKmC/IgBykOs98XY939WWzIPKKaVK34lmZSIiU35fxiYsz66r95s9ZQFy+vfywk/Y
B+2UYbxQfpXW8c3mqr8l3UBfn2DFFMKWBBLEAS1+RaP1nkiaS9fTzUv+uwyzJVg0jNEnGuxSM3oB
l7BbfpdhWCpfym8GYPIzqj4gDuAkcvILfclOhJvvnG3tOeXJsrMLzpvA6tixVL7rdZMqjCfCqPCP
SBVCgJmSPgS5NxYO8T0bFgZ1E1DAPG/pjpOg5uo/4i3EErqqQ1tCdvn+1sBz7BP2lZoM83LyGB5g
iItYr9TCxigE0SdkYY5+lP93nFDCNTwboYu6EDTYwnjy+yW61Ih4H17/TMg+vOdGv4g/1PdtNxXX
5XGCX2dG6bTsKeZ4VswrpiRUjJV9KGA4V6yxL6dZI1KJXpxAsL7cbPrlCCpoy8BQ8Dpjt122BBzf
fmAxI/n1fQbI5U7wYxaK2MzDrFbI8ShhbeHmgsCvUPWIubWxvL/78MZYry7xcf9fxylrnBl9IoSq
TDbfDbDHww4pSBz/Gpx7WvcLBCk3pgtYeDdBd+zRvH/QFPE49kdx8gKnLeyA8TxXFg7KAMbNwgzm
qNjNT60aLoxMsthgCPnWqADzETJWpC74VOw9hgkplIaryJnMHcsXfCArwmib+t79ubP06mxMFYpH
IQ2PziC/KlYdRiQ1EIc0Vr3twD+c0UxVKMPZjefBwZzyfUHIOV3DNAeC2A9J/wFO5/8PawwxC8cG
QRgQnhU9WWGOg4EWFMHktgY5r21Vx3Gam31cGA9znIWkGnlWtcw/iQSftZx6T4IZonkkPMhgrQ7r
Y4XMHrZa9Try8WxCrdmbS63sx1Y459WU2Q19XfQI9qSWtgqzqCAj6ZhSLz+N0DY8wVBxxath97hz
OJn2+2kFhvVLdPcTLgqpc6pMLjAq3pSGT6tllKmBoCA3+rVBVsRFtf4ZgWIYdTM7YTk2Y9olgwOk
VIck2qlx2eRlTZvnw1I7j9DHJS4IuMHm6qM9y3cTSABIM5YhjeDcuGjVroQDjrtuLuS2D87cykeF
EhQvyl1py23xl/e2cxlhIdaPl0s+3j9ig1t0vPp/012YvUXjCkoZxM62m0g8mOOGlhnCVX0Z96zu
I7vi0rQUfRubbTB4CTTphjTAngEN1HvaVgSso9sT28DMeqba50jJL1ccuRTNdytLpUfX5He0HAIW
xwYLhmR3nxclSifgSqphY6DRb5VPjvGIHvcuev3GEbHjSdmHt1YdTGZOknOvfz8QJ23kFBCfrP5a
/noUxjR8t/KV9YQjuGV0BhynwgqcNjYnFYU26qnwvyDaGKcFqn5VDudMgYtXxbZEKmVsIVnVO9D5
NBY3Je/9A9SZEVCJGUJ6DTDXB09XspaxeDXQmIfkEZmuTGmd6PCydrX69UvxIRQClQD11wNNK8xy
BGy3Mtb1jaT+8Dm0vlIgy3cYDW8s9S2a39jOkqqvYh3Sfzw46dn87ve6Mwy6L3euOAA3O/FqwUOs
a8vMQYiDIePvSCcTyZkrUcNVqAY9RZ6wENOH3ZhwUB7AORRrDXSvcyHUpEgEDecRxsZ2PogHS+ZV
AhxsuBPY3jcOhpaAkISCHVDWbWKPYWCPJUZqAMeTZj9Umy76bg4EJQ9+76APPjiupuHyuYWr34pB
9han2/I6M/YECY0J2yWvzQHYTAqfmwEmoZ0jFufijxFBLemn3v9R0j+n+Cug0nyXEJLPn1tCStgX
dcMlZGbvCA+rQGPZJQYuB1Nabc/vmtdUbQ2P2b91Knimm2yzyPw/xvw223s8NP48jiD7uaAgB2v/
wB4zk+QN6LxpLe3+eNYX6BuY4sIIMb0FkeOIZXfvUBxvZOJLl8DtrOBj3jdp2gGdxBu5oX6MPzXR
FS1GBEcC9kRgLNl7yLGf4eNip/GusK0LiRFsR0a8SmzpogCFnZHQ/YfxfRJ19C3TMzRis5SeLzfE
0l6Xw+IBCt4qz1HgI348NuF/E8HzlAxA1V691W5dLBCMFvh43MuBxG074HFxKyJpfNGXcMKwFuRh
ZACrL9hBnARnFa72TXKhVRkQfwP81HxLTo3MC+OBt99wSYVeM1qXIFTnERjhnjA9oJC/xN18lYmW
Wx8T9SPoRB8KnDTPekDxCph0nPQDs2nJrn5YnLQpmGom0WTNBLpMmqvQprxiBmDLHtxX8aNHs424
vfnpffGNnyuesyXKsS8zrOGxcveljkKY2rNOgof1YGA1sUCjNz7lw1p1XPv03xbf98T98RwT98vt
c89U1lVMDGNLErn734vS9/VjJvzEZ1gYC3SW8r6yLah0vFu54vkDMCQy3ATegWzyoKdN4Z2JvYtg
9dy3xiQ6Bu7FQaEm/kR1iUTvetq27NazNQTpxYUeeNh/qX/29VlSB1jACfrtGhQ8U94rnoNg8e9T
vjpzUft5qLdyZoGrzjcL3w0Lubif5MTqKSavdtQijVUTTB0ZqLG2Ent/dDzgOndI3gXbl0cWvH7Z
bj+CEVowq3sk8UoSF64kvUuVPi8vt3qlu2i1cHPs4D9EsYTtWwh4ptzKUVGnVn8hslxJCG0/YLUD
fE/plD0AV2i+ieDMqxEHaaY2dHHRnpyePPqlnNz7+CKa2eiJOyks7WXzW1XbugoumHsfZi/GOxgL
4b9YYgNVh3HDRL0m4P7faYRI5nwQQz2sLHOyUO56Axsw3shz0D2jaPL6uch7PP9BWxeqZiXJCZAI
o5U2TeB92tpVhE2PFkCraW08l1UsFABGhVVMigZVHjbkHZ4U4Kw3cr7wLLAZgf5Hme0V5Ic3y+Fn
WBF6MwLMOB5mx4sG7Ri3lKKS1TFMBA0s1lfR2K89fYSl/WAJI/508zvb4vlVbNUbG+TTekJQSR8U
1LAffiGWIT02DYJXAXuaDzr3Fy8Vg1qbGA7YUjqh0kgwVulqTjahMi0/sl/C7q7jVfbkxqGSze7q
wKCAMCdJUxnBy07gOe6h49gBTXjwRTmnU+hlDBSKkGcTlLFHHnGPK6RNBfhUdvqr3TAHFhPpZzZW
gpeUqCL6adrzxdpqpY50a2P1S7MGQ1m9fqYldsd0/dBsNh1GL4DLerWTI6nF5ZZx4EzSpK4p2JIM
tYwtoLtQoLYg9HF2scUoBViSqawbtX/Etu6PrIYDn1L9b9bC5Avir9L87/6VEeHwhVH0i27gJtX+
yWAqfgYlDSv5HCYV1bXkMkldh/vS+tRFlEUbL9HkB5kSClnEYg/pfrsieKuCgR6sTdQAtK0TJCjc
DYjbfMrvzNDOM8xUAEkXx3t4svEyudHtSo97rEA6JQk2rOU7mIWH6J4yTTiYcL2fjMByOeXFKgOT
BuqQogQ1ZgyQlkzqnIeoEQvzaCQl1iZpkC502M8byShsPuPXbJYOvJ+IuW3lMfAkaGrB5Be3NIBL
iFQCvaMK0qivcNnFusUS/IUbpzluCSz1D7qQ3sQEk0WDJBySkqOVnPd85gER6LI+E7XKmcQ/9+U4
T0B1k3/clfJW3Eqm7hYwi4hvRIh1awLxzJwCOzu0z1GKc7GBl37hlljHAZMtsWCwGxEvbsPwS1Rq
ISztPbFi1q5Nqh7BkkrSjOkiHF3TTcNls5Pgk4ZV5CPOzNNYhVaoUZf2u08ZOGfG7iJGVg1S7UF+
oTCn2NR0BrgRrDS+rhmM31dyOD33Cjs52wX/D85K6/m1HbY2iVhz3YgLnFoOTg6GW+OQnhyOy9gw
iOx3SWISh/3CCJL/vJosKZv7diKbPo8PlBX/CGThr8zJeiSvRWBTCKQm14na+8I8wGUm2iIbg/yU
0UwEamP8vBk++12LsYEv559q53zng/emfThCQkygwDp94dQdh+spc1qeajSEFZKSQv0xVZHLd9r6
3G12ec1XvGfTmirsJkZzdLJC2fr/HWcNrhZE7rdcvGPqQLyktKglj5rKekSblNeP2MyVM9Okc3Si
F2aRJoth2l1g3Dh5SWYtDMgcyQOhXl5Nj2Xr+GcVkhZyq7QsILQrjytPQEWUYWPR9DSX1AvP6LS7
hJ6KKZb2Oq3Mh5oZOEFLki/ra1J0ONodhpRwObSq8o/KD9nAM9K8CHxD5I4+qdItINKpkcrbQYj+
eXVJz1NZbHbICfs8x8EhiSQar8g6WkfWP4LGhOl2mXZhVDjvR4NF/kMQevSr9Kc3fE2LjYCqclF6
a9zqkBfIYLphv1ehyfX2HRmu4gMOJj1cwIubwliYLB0PvboVJgHgGAGUU2lbxYrFQfN4NuOXtj9J
AqTQE3gMsoKGVoEibyRr/B1XLtKhLcdRkcDWSnMxQirEAo7Bg/ba0ep25lCMqWtizpcbOrr9J5x8
314wcqh5Z9a85YKqrXrh/4cXZ5q1ZWnXIInydvUhu6ivFiZqQsm6CkqnWVgi6eixWB1liBbKxxXB
/hFgcoaK5vu8dgDcKWJS46ALUby5uPr+CFBI8/NxGXrvPhwKHOxhuuPXJN3EVMdduG5/JVRR3WEk
Ib7YX3OkT09P+zn0d08NUALeMhNX1ortDKPELwDOGE8Rl/AL1AOZr35CdVyaF2nFjhHnkDrVxYLW
1nA5+Z/tuF9U4YutjhDvlBY3gP2tMU+Q/X96lpuQZSfNlAPNjR+tl91C6XgkaNfXRiXH8mL+A1D9
vqJytDGXoEa7bVkHOc4JUPNBmzW7zUfkUTtP0LSyL5PFPNk1INKoD6lqUnCkYBqxgQ+98Oj0781i
EFY6dvRxU0S2e82rvXXlE80nL2ZQC7IeRqIbeYZZBb9xUuFs+7j2p6IMyp6yVfbykz9Qvt6uEqWK
6jiq3nGZKrwWjObR5IZTfrj2jNN/DNHbJcg4ljMMYgda0geXGkz6nK7KM6TyTwjrMFVFpbBdy5AK
Cv9gHbTskIG6aV5Sto4PQY0QjMgUAPISb5taCWEKf7GuSrA3++cElEsZ83ONTOCcsCLvtDM66dM/
N9Mf8XGU1rZR8WgH0utmhO3bZ6DR5iG0zKNJwxO8oCxWWdvdr19vNgfk4tP6fXoLKJW7YLC10gY2
Cj+MZDDJI5xVKHdUf7rY9i8hTcSt6a+p8lJ0dnkg0VOo0BkTkUyAKK6M15sl25ftTUHTx2lG+UG8
br0B9Wj9nFNXta7Gn7Myc/QeQGQztvUoNMoNgeWXNVGhQi0I4UMjM1km/sbhQz0hF9LyEZLckPZO
pHdfsZXRFkuryeDN69VVOnoOtFPW2adyjKWbOl0db/vm++P+v9FXLgs+sG0qlb6gowOE72lD79Hg
vO3goibrvseQjp3v5crocyKzc9JcdD/3wn4STHAuUzVdxuSl7QJhkZm5UYG1O2MFIAv0W5N5v4/7
Cfy83KpSxayGpcKR6Zv4yt2nfFGCv0Rwh5Ny1yBpgrnklJ8rDhYw2X6TwnotY41N29gkEUMbSiE6
Fjagi/UZeDIiosMhTz74R5wAt5qNfMtnLFRKxRP8J+IXrT74uivLgEvv8TkBE0V4ZmVuaqLNxaQO
AL017UljzkwvNiOBO36il+7exvRTZqUj8E5xCWlo3zqrfHZLJUP1VjqS5ORm/DZvqW0TPxsrAY+K
gKKssBb4JGMom9YPVDQpcxrI/x8Ul4McMlp2DamKWeqeq4rha4D53euj1udKXCb7unU5P2cuXIxE
3IpB9BA4ldXvW1pl4lwnTOYtHMJ8xxDmx8JhfzCjwAGv0Pp3+6Pf5SBW2mDxC6trBR7mufC8DLbH
4SansxsIz/FvNXfGO8vUUWvgE6iVLbARzt4MwhQx/knqxRsvM4/cY771emI5jP8M1EZbznt7PzLs
l4N1tZcgk+EYcVe0NTf/jWcStjsWV4Sao/p7tTa9dgO4UpuApF/MClEXiilog5STzITuZOW1YQi2
bfo5BuZKg/3osL3v2tL4+miHj1q8P+KhEIFnKEOP2kI8EOC35hQtU8ivAZR8mzPnshYG+TjJDnc4
EwMl8a1Pa+MqV7Q9n4MuUgogU4LgtR3NT+UtQWNagSRRGzGHgLUPJZeF3r8TUUCWkMeFllvtSuq/
LHHiP7CQjO7SbUfh99kzb96t1WA/suEcNPP4ZmRcn+P0E/2UIbENOhc/dhZnaqaFKUBxDcZdR6B/
2K5d7K3RLkEJZ7kARz2uHCUF1p0+raStdWuPpvt6NFDjmDHsiUddmvpmQo4Njjn3AkPjrlXF/wAg
hkQh5YBHXYyMuHw1DPfMOBub9IZUShjI6I9RGC9yFwmePVykhYyxwzL6nREi7/DX+d5imXIyFvdw
R492CoJ0HXPiXgickDaO0b6IOEc0HUxdCnlOMkk8zHa6kF+a4W7Cz+IVydLUNoe00gmW05/yIyyD
60FQGfPuEwNvVb2yhhzrbZ6p1vdFSo0UBxMYbNmODGRcUaJ844OM/Vt1ley9/8GZZ1hfqFNTTMsx
EqGcP5kDGz7VxyRLfMNcO97qO1CJZKaLzFqBhQw5ZUdhstT6HPiJ7a/hszUMfVVRsndQ17MQwZUl
voAzySaqyJP3cQzFXkdHJxRvuHzelRAzvzJlqE/f80hIi7skkknDOpJILf4wg30GRI7kBN68tAww
ssGMVtawiFkjYz2zBp2NLlTeMi4fLtAs7qrJccro+pvOnW0vBgcquSR48iKRmdJqlrbXpHXRl5In
CuifLJcPntaANtTkqCAg5lB3O1gnlS6B1gcfIk80Wv/1II9qhPYGNP0dnlsZvWVw8c++ngkY37AG
XzluIO6zKeO8sFLWpyPDhbgMukBRdbTdE2PBcRajhhQK2N3+Vea/gnVslQog8V2hh7ZH+8hTIjRP
HMsGH5lRrv8sTmHbwHN4ukUfhSwk59bfW/cU268Wy90ONIbh+E4Drm6Q3AEgydtWWOk0LhU3wx6I
TvLepINt9btrAMfPq+hNSweYpjhEEVImtwcqFt7c4jg4eaj+mOYfZRd1UPn24hZV1Fn9yBNAnX7K
s1DJlS548pd/LfqLJ7HO0I/Ai2kIUFV8KJ+ZOBPy2t+HA+2aIGjYSbDlB+aHVhDCQg3F7IdUZlib
E25us76brgeI7Tt0U4zG2vEtFgBNAUKDfvZhjPyM1k5PV6QPg1vqQXFBzVyWT6WpJCHl+k3Q//Ez
QhdALy/txvBV7Foz8PQzLzmXSkyXG7rLd4PORag1CsFi7Q/1HS8FipdUJfVluj8R1HNiK+bfhkTF
jw11ASmWWxsDGvZTdE+2i96E6PQQgfDhpznCNeEvUGKohwHmO/rsuLv5/BlW8CCWCwpA2xjz2FAy
CdW9u0BN6Z8cxuwYUHzOwdYLIRNCKG+zoGj08DwBo0oZvsq5oayod1EfPdegg4vSX7YDQPExCyUR
pztKrn3iFEYwHtnbevm6X01couLMn0DD1SnMXxmbxZjdmlBkpCLWBToq0Hk3n3Tp8TCo+wa6Iys8
IfMifEFm8SQa1JVlYbuc+AqRSria+igeMMo76lsODLL7Fapc2HYgm3RewRU3wUKN2LZ673aDHNM5
hWo9NYHS4jumjjTRJWgIV9pI1SJC/X2sQLnhRPrJgwviM7YBDE7q5MQeLqUeD9dZWjVRUzS5VDNl
ODMUl/LAO2qUbwhngIMrJPTRjNYvZm5d3bjww092A44ALLrgvGXLCwGqpQTIZkHB6xw3g0RTOULp
W5nhQa2g7wcBGR9p/F3j1EvsA7PONdgdm3COriovOnzcpdDL8Y5TYGad+FmhEE9bqnxX54xiqY/L
Htoz9661TpyivirEuM0g6Qog8kFJCl97VrzgXKTAb72Yu9fJqn2mVEcA7JRmwl88oYsDhL2cReWd
HsSlr1emW2PUtTxQXBRYwB0KGkxJaKS9t+Z+IEpLWd8mrmawXz0eXXkDHn9xypg4IAMmudEBao2M
M761DWIroQ1OqhmoGgGlVzMYocxluI8S2uOyQAGbyKB48HuuvqIkVLP9Qul7TbUoyvHm09amRueh
5BlI0UsF8AHfVwolDU5KbL0U0wmlggiL/PnP5M5rPm6uMeTmW0zjZG8mAodgzNEuWCUPZYFkN/xg
EcLoNPXREZImAzILhdEN4fH46vYdRpOPt+iyozk+4R+JVvgL6+xJzlC0eohvXSg1wEP7xTNh8gf3
Vyk17LvPWM0jRkt+VfClOlkCQFoawArGrYjYrWYh5/+NxgEgiSgIPKaolXBijj5+Budk/VgOQe1d
KTAGHgCNyX2CQocDIPYNVgRcSzVmIlNL+0nN5MLGUNGFAkI8P4QW7AtJw2WEJPDyuZ+uljzl8lWU
eoh9lkWHL30H37w6jT3WV2gJf70ipZhN+mVzd7bHqNQNq79C6FY8ZQjfsSuEm1s5mA/tt221TccB
S+lndVMXUKckX0ngrFjJqd2Jnivo+Bchq4G0pd8C6hnB7+SmKuyUsa4qK9+2uvupza4DX4YJeGe1
TX8ZWfsZSVgk+jqtF3ZfMMYw91VBKlVPve64f6m0yJLufyN+oMhqGztKakspzZy3YVYlQAhnZI0c
ogk6StTXv+RCPdOLoGrstGRwVDElKMw7UygnEPVeOncvqW0Z0/ApdSzn5AZ6CniFGPfsUisiReEr
AvlQNqdsJTORyrtj9MiVP7ekWvOp62lEopuQCXvt5qZPmVr91UKEXWaCaIrsj2KLbvSPjTf/0y8Y
a4uK1dS6058e6Jpg9ZtvHGgv4rm75YtSiBBqEqUjotTS2PwgrZI1wQovGP6t6x1V51Qau2SgaDtu
vT/ROy0fV2ND1WiZvDx6FcnOX5qdvDLznIixSlqwfEm40mih8wt8KAPFWHmAwc9IFsxhPXdBLgQw
2OQSp/EztVxNfZXZ025HLbNfMz6+gTGnPKBvgj5YcZc7BOalhZ75rFEeej1TVaOnfD99JVi8DsqJ
njRTAP84Eir1Cet/6EziMi85CseLeV5Isi4/hkRnid8OTPvZjs9nIEbQ1lIwS9guqa3qhb05+ozF
Uh2E/Qp01c/l2iK5WkGxMZWDzdLjvb13PkpDgpjlplTBOsUylbKGySqadMgUUbN2kcOTiMDD58ED
p7+MTUwYXpPZYCs6EX80f6l/DTM+cxgdDEpSI6DeCtYdDhiwnyRSqXjTAaUW6nzvwuqiRGIvGi98
fQ5RAFpKrKC2ChjVJp3Be+0zSyUYi8ULjK/5dCKKT3a3HXfdFWYKwxsG3P+8gqw9CjKC65TQP186
yXtt9iTfcDlCUVFlfJqKuucOhHoaKdgmIf718bRg4uXwwDWAgerCZMT/iEZEp12pxVlLy2R949Pl
AoDv29poYxDFt8sSorhTUV4+fjTa7gD9awgpN7b96dBTyhGHbgkiboiMuZAoxS9tTGO4WtaeMuyE
6AkGBujHhn8SzfdqpjQV7Vuv14lMRcdh4aysdAXxltPgqKHWDgi0gW70dCo6m0e3ai46TiVB0pwq
7H9N6rojMM8yq8E0hDB0xxXIm06x9K2XttAq/7vvxA4+7ejUosmAYZsFhhsYdYYJMQJRYJjsCvu8
Misv3nWls/1+lsWYVogL/kPe9gGv1J1V8F0UhK1h9m8wsK9g73fj1ppDEPDnhs59jXzGzVAEc6fQ
MiETsq72Bsg3ETQWAkbCixzvH2pEDSI4tVoMfCSoqkW44hcMsx3suZ0suelfmXF/z53kxT5khJlp
M4h10zGCgO6R6h14KB2iAtjf94pmC9taeIgoaIJAraUlSvPaNeT+qQMg644HMmmLuyOhHY9f+duE
ziUa71m7PkPJcGhk1nfY0lj2XMOkB1fHfvgo7q/oCWZ32Yu2MjaU+5BZp3xmst+jqj+KZmog72oM
7Aga7RuqTC9TWaJKjBTeURh9qCZM7WfSawxfPqli7Uypra0q0eLDvQITRGXc849zp9XgTRyUEEYd
vcuuHQG8Am25AyLCcgwZ4JCyqRzF28bZ9d0VvYOOsh/5dDVx2jdESoYKxUaYfgBQPUdsbDNNw1UP
dCw4k869+SI2GtqRKnP1FaF8kyvi9YiwmRbeKEmcIM9fMTHbJENqclVuWalDMoLglyzZ0jb0aFTs
hnFTj8695ysS8OdDSj2n4B0YvDeuwFu++xzAKyyia2utUQriTzQCVXxNPYkvlzLtNYhsBVJhadui
6UlyKlzYu0fkMXP4xcNEnLji44y4MEqqnerh//Y+Lv0OMxk2mjOAGJqXIC3X5UAAssnZSJ+T9GYi
SxcQJaNH4w+wOMYsh0mQuIOSwQi+q1fvM+9mWOgEDYgldKd2QcT+qEurIFaf9BOsVAl/QJKtqgsr
KDrm0EKwpO4MGDUcn8wxdqvOSqq3WkWbHKBn6U8W+MAIp19Paii1gzM7T9Bl4ScODZQZ/559vw2L
twgfh3Q1se7K9XwViOMnaXiq46VXNDYyN3mXXk7CGMx/BLJg7Rhbqdbs7qSyOtw6+Nm+FtSwGWCO
G/aB4KKwQnND64Xj+ordkCPESIXHLyX67MWeKkG5E+7e6qNsDg1zKnr5YUNOmzilRlCS7znvIAnm
Gu1InqylpMOvnl4ycInXb+m+HQiKpdT1Vn7TdWF6sUe/k5rCFAJB9kmeeePwFXdKVLw0Mbri03Et
HSApxbpYZxD767xUheJzewzaRTexldaPhAzMcT+K526+rookwER6zYuu0PBpsSIAboQyXRTpXK3J
0mnWMNGKTkOQ1jUvCnQHtJAN5vwDpDeD1sRNKQ3LXkbRjJSkkbesc5QGS8G5qHLZ4uORqBjQX1LU
7YoljDhQ+ZUxpSiHcb+mLcQi2tyb0LwQwdbov3pxnqJcBoTw2UkDusJ/oNQH4/iTYcWFf4jgUTBK
DSn/puamtxLyqcHigcjkIBntAv4PIpn3E3VWgRfMN0wU6l1Y89P4sNtLatc/yOd5Mn6nwuWkVt1R
5fAKFWjOtOdXU+lJVbjUaA6I4r8Y5GEURmwDCphr/YmrHZGttCklsuoHsexMrM3820kySyeFoXDp
s1nNq8+SKrOYuuvhJCSh/p6O06Hx+2Y1YlRmueUHiHUP7ekKQVEqcSgsJvIwFoVku7ZVAXf4+e48
ntWR8UAyGnLiQcJLd9IcfiWGE47cQ5w9EkReYpl4FW2mhaMZ3s917gDp2vQNnT+l3JM1haG2wVvX
SsdQP9ogSi8YYiz0RocUgYjkOZb1aAgDBTHQtjwSTJPr8ly2clXEitIhlVlGlcFJJWiNiaXQfL7X
a4AKfvPHnFsS1P1qn6q9Yi/b/s5igkltKadcf92tJn+ax8yyVQPtniI8N9HUW3AyfaVGpniUje4l
U3iPJ6lE0epSykjuoB2+H5iQRZvxqfQW9J6SAnrDYhiMILPw6YqWtUpg4cNsP97bh50gru62MF0U
rZA4notYJYLDMToOkhMqI10NiUnVmaiIeZk5bPN8ah1Ip09LP+uLqqGeQCn0g1M6PsjHCgavtipj
zei4n+COBitWpz543WqPM3vUC8BltZq242p+buNDxwi8n0gvvsPxi4jfsPsb5bdPSXXGoAegG6Nk
oH4H3eauZw0BczkdrybDv+SGtvDrhYg4Llhd6+0RqKXHJNoVV9Xg40GJ9vbwAreEXI4iB+RjHAJY
6Fn7W6mAtDODx25X9yS7iaKScmPGE70LvAgN64bMQMfOlG4oKqq7OnuIcU+l10zgbdSQaAKtx+eu
Z77QaOUGbd27dY+6IYBD3Gk/e0sGlY72Bf03dxYYYZvbZR3XzDR6rVf/Kz38Y3cNSs9UNIpRndY/
3+LDLHAzWj3PIiRiBY56RXoe5JRBs8U0qy3yYiTxuDSzZp6OBmW+TUfi7d/iCyYnO30l/HwN2Ety
oVZ3iCtMN4rhzPrZ7I9p8N33APRAMWcIWuCdrxhPyy3YaZVn8u4bj0VnOjivkRlpt+EdsZ7diaJj
80y29at7ON7vRb/y0XckLlj3qrTEj7fm1D8CXlQkxA5AFpvT9sqcJhlQ1LK0bgH525Xagn47vzWQ
ufcX+X3NqiHIGf7XBuNVOoQKPs/E31VY6f9EUqZY4Lx7lSBSKjxFjBsKzVlDCAgGPC6t0e+aUyZd
qBsjJ/4HVQOupaenVy3dhJb8ShIPb6618z+Lkvmibj4bjNCZzPYUN0Z1QLRgxqtFpLGpOTULFi/Q
Mk+JjN9msoUiS2V411d25nKSqzDO/ThJayRQ6Bc1U2Qm8miJcrgJ87APBljuaGGRwSZB+WyiulK/
GUPgDiyTiwf5rBDPIPES8mfKJy7Wn3FKQfcs1+eZuoz92EWQwLvNCHeweo8YtXt4qNbrUbFavmGQ
J9/r4UGAhziwkX++GYMG9URjTwN8NUh0vzWPXXJq+X/Gn10L8VuMqBEOw1PJGfHUfMGVlf8xbox4
vW6mSlyV32VVqKgS9Fqj2RR3oIu580YuSjUskQfvoYumKJNFJfz8uh+vG3ho41MHWgjb00E+TWQz
mnkQKFwBJ87J6yhs9/nY+MNZAyKE8aZiFvZQ5L7S+5yxBAg8VKhMAieK+fYUfRzQG0mmuXOgPASG
n0QXaYzvDjZ9ouoL2+tU6Ac8Xu5ZiwRAjrv3Ct/HLbH+owZEPwHr8yxngN/qSmBcX6D0rVbMME8V
/ey/G+JouuHWt9JAlUHSa5pcUZJviC3iN9NJnj2CeRA3WkcY0TSEqxAh0JOaj2ELBgfqC3vlkm+G
2rR5+l0zJ3S5gq3jjhCw14MRr5Y7chZwcIhZo1oyw5xaxPN/d37ByNKGmeuIDmqPu1I3tVhHI4h6
6eAyhzFDqX1XrxHRPJSzlTNxS2aLDXjYPnL6Kg6JZ8dGMnpqJ92GMK30UTb5lunjHWzY0e5fDxgT
Naw1kI8ylFqntNdZk6Khm4RYy7yU/r3srnMihNZyka9lTEd6HVB2/WqdoB+8
`protect end_protected
