`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mJ4XLEqtCDcrMYTrTFI/GxYlB2EmzF1NcxKlXtSU476Dr03CXhRO5LpPp0YK58yuwxszuRRhfcbC
tOvm5I9vmA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D1G+VJ0wJbZ6WECZVA3gAfjyRlinciGD6Rv6LLAAljxDndve1cBeRyunJmmYLLboRnbqCtmCTy8B
fWff1iu61CQQMNb4VUoGG5wl3q956/8TQOKQXdCwdnXF2mS4IqAllBO1nF4fHUltbwzDLkmPQsno
7eOBrvexQBCCSXrznXs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
COaN8aHyP1h59D+dw/Mr2FUCSZkr9txgX3aVfQw7BSruEzvAujunBOr0qlQbxnnkI/zCHAk4IzfO
Q+urbjbvzLZhJg+W1zfWDMuihNJ3kMC4EF4MPJDA5TNhViayG2WvsuguksmozCKYBHlS//nx/Wd3
LD7K4c+eo9Xq2P30DPEo3lURDQbl/+/NfZloDLq1p8Gk4Z21Bgn9b/NfJgCQXk1839PvqQQxi64c
vGcuuUDUg7s8rYAl9NknaBidpY52tOZav16CsVZIVNo/LpUImTpIhxZZMs07/8fjvR1NfxJfQyeC
EHP30jWxFEfN2olQ2H5poOoRgkITP2GnbdnKZA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U4Xs9EjSo+rjqcBj90EOQnGF9BzuGv2ZMp+3gglubDIBbSoUej01z6CCohjMRMars3w6GBUUO5qn
xe2StzYl5Op2eeiqITgtqcGcpRBNUVgzFyUQU1mr1Uzm98uuSHNFjwndwomeA4BcAc8c9M/ANIew
7I3QW4yF0wdWPOUtqUA=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RlaQ72WtqEIOQriI0zYDRsxO4rBq6ACjJZ+lxozX7EFWMWyTtmB8+d9vAWcrWW2Z2cUrPSEEv50y
go1WsufzheGm6JRM/ZHbzcerQ7oJOvhPnDrT0inoseLFEhOac+9X5eZZMJ+Am1eTdiRWt/GhKzZR
Sftiaom/8/rALYXYR3QK/9RaxfpoHLGeZsqYlRQy0NdXMvXhqz9sTtkBLU2O7bunjf57fFjwl2J3
EIhWxZ6b74bUFmu+5QwWSBsB32NXx4XJh5B55QAG00e+5Dr796LANFrU9UeihXH4CrDgOOj4Tig8
Cf19fNacyC1UcpXrgXR2i48E2LyIPRVTzjixLw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10112)
`protect data_block
WtaZQ9iF2AYYrIHuZ2+RYF83FGW+DGnPt6FxbL8iqao8MzmLem6iP14fWyTCjoUll7qzfgGV4UV3
9mwkVwdXdeT1dKfprAKLbA1yDfS8BAkFDTAMmbr6VuSX7HiolL7hO9kgJFoC5AoJX6oJDQGqXh4t
qCTBbY5Z6Y5Nj8GHJFpjHsI9AN2CEnBmVvwIrWfR4vHWdNfihVWfVjy6K2LCzaPyx1mNDxSJiiKl
GH34DLmtusnAw81ZmxzbYmUfqnZwBq4TJvIS+PUXPORzTH2a6xi7JfkJNwdXluvQZcw6g9c5KAlZ
xlRzHw6Hs+YQpTbmUdWBsq4W1F4RgWcS3H3KEhzGPTRqkWzJZ4sE/LBEPkaWKHCnEIMw4Mn7Tv9c
hOhytwcw3vuhd/QRgJHcG0MGY9NUq5s3y8naV5WQklU6PvVJasD6LcKsBI3EXG8LIFliVusmVAUk
cefCMhgfvnqzERQG2qRpcaowP6hrJoh2ChT90ggtJxEsKX2D5jyriKvlY14Ie0JuM3JoujVmiT8g
G63cQXHKqaSpe2YwSmJPRD6GHF3VfL52wwKfIWim2gOwF/sFkshVPCslLqE7RXc8+cU4eBDKsdjs
uRmNrErDz81R4POSazC+RtiILN0nCZCsobCaCRMIJnqsFXVs5SH1fOohlOoEyrD5cqnpYBnG0RKP
YPj4fuhvr24O0vxiLBvQKwW/MF2+oMZfoMWNnvhfauwElmw6kAI4jiTe6lCwt+uiKd9uIu/V70l7
/buHVsHSXUjm5DjBhlblR1NNVa9dPAM5IBl6FLz3hM+izfFRIF2et+aw/pTKaL9hfYN13TAELdS6
x3KLx3mE4FSHZ+1CuQLOK5bYNeDB3qbHn7UYghSqGf0o7VeAm1MAcGfMWjtCpQ7crR4UBhD8QS+d
pNykgSM2ohcNJRXHQ+Jocuw7Ac7pSt+muy+k2uaknXEeFC7U+6lPT2LsRQjJwIrfxRnPhYEj1KGB
MaQ/+S4dIj0e+LrAE4MNAKCMr6XQpy//GBM0DSK9RnWaip8Ap5cbmlOSON71z8R9Nr2Jf4YtE9dT
eQ7Pj5gAorKu+YfQXZvq2t35XGtnVglEYWEClktWI8o7n/0jcBriwBuGK5dn+l+O5UL9QYK1Jxv1
Fj7sAhpWeu9sIerWMKZ3NG43etAKOXNSO+34N3kB/RlwoNEPF31EyBWf1qkwCHqUahiRMKS7bDSR
I6YBwZOH1ScO6igov0v0vdonubKSCp/tpF1t8MSegdJSzM0G1PzwJ8FwVkgqSRRxzgFKYdwBVmUI
2+9vvAikrxs+CoZZE9NrtzrHeGspzy31g+zbminlsykTsSsVuhKVjSKilo1jjtMAxpwJcYcbdqR7
HE4Ihe/jNfUiIxnTtFL5q2ym/etb3uj7Azg4/lsHomVmUx9hHxkwnAyXx+UtMJCjo1yCJuYDiMaZ
NLTwV7uEnKMFdgvAYU+Ew7swTrITg3va/IsIL992KX79TN69DMO3do3xEQHQKKVFC6Uav7Q6fz2Z
lb7qyxwP8q6jm6WSu0NCyja2XiB8LIrsDXZh+Qy469xUt15MHja6wdrDguk1uBdcTBq1DHGYpuGf
xt6PYJd1tL3Nnxag6YqyVivcUeyJwzqd2MYzfQRyhLiDPmFHe27A+4GZEX2iJexK53lfvFewtFWe
n1PF9nRQ/+Kceelz44qpIlE3d5eCsPLq/c1LduJHPw3ASg9xepkA0QKrJ5X/lnR3OGgcOkxY4FAl
fYlvgSTlcCSH+TxxFmngyourZ88KPQCYUc1UKDAA+OJkrP/UMW4PGhYViY897hawhssc+J/lKkp2
jIvb7LLLbLrDIpWTbb5yxN9ClwRuYQGAf4yxHM6/m7UU1ChLaZk4pLMtV7K+QpRH4mNzPXAsvSb1
WY0VkOHWaruocq16vvfCTWVwlrBUdB+nGJjbAQmXWwxT8HjSnxRGnsEHSpIsTDulnVBf9zqGjEl/
6TnxRptBK6VCrlm2lKtiPRX4rP7m/0e8kIg4d8fqNUDxCvdooQF+p4Qi34hMHrInG1IENyChiF+S
L0K+Yfre943hLic1N2/rlDTmIQ7B5W28Q3kT2JBCq++HGqUbuO1wf/M1rubIpjumgZqoQjspqVNU
6NJKpdYty05GjrXEOBjlyqELJo71/L4o1yhl9paPUyaBLiY2SfbL6Ba6f76U3elAZ84LJ9WJkRQP
EB4zm1TiRDuZWhF+ZRsxXxHc5nQR5WOZi0QnIy07PSHH1IvbF9Rw4/XJni1LNh0JdUgSkkBfzZxB
tWxi8mTDY/lHzk/99AtHhKN/+gPP0eySe9G3rNWRemLqLLguZ9BIRreeFupIzgnJNQJniQzPvZ4Y
W/fEpKW9XSLxHwgbEfSU1xks92aNfl4rwrDEyj4I0WLeekUxd23vc+IbTWKAl2lJgz0tbECnpDNA
gpLlMERCwFvN1rOgb/EQUrKtY+U3JEFdxNyE8GLk7AIWzO0UCuoVn2sz12ilPY2sHUdcUQyQc1Cg
tyMUPYfs/lJDguxG1xtaN2dKtoXVUg26fPsalWFeHgIDQO7cV0X0KMYjz8TQ6DsR7twVF4SAshj2
z4MprHt17pgHTlkbhQsVXcexBug9nbBtltV7dNoYtcvJa3acrKg4pR+iiqvm+oAdstcPsCGDc+Ra
eC6+nmsvR4GUH8rTHfLMtgvNBSWy3/Fjmc/9Kaetl+TzQUiYm1QhAiUbnLzVouD/pxf7jjpa1gTo
rgWPR/FMQBQK/lEwy5UFXbE2tTs8udQM5elvimvE3aFfGudNcygRwLixUCRewIm33DNAUyC60+N7
x62nWWCLmUGaY4SWIqBbujysBnNx0gezNZFXXSTf6QbpBSGaE9jBX+hB8C9qJzhBWDAZA+8frmrE
mnJkVpsT9rJlMAovR3eC3/2bnIL6Nw10J7/3uTgRDcMIjCWL8T7I0fR1ayBBoU/5kMKWnaayAmtM
kO5fO9PogCYd+D6kVvz8Rkvyf5ifAuVRCBEu6OvRlPeKsdN+V4biB1Z9uRsnR3kUl0V2tbND7wIZ
SD8foQZny6dwIiVjVBy1bIicF7MTEyV+vlQQfyQ2BoMK/0grq0FI+5loMkCn0cTWE/Xgi8ehRo6C
zXMMUDj48/mWuddah9Z+uwYRhKpEqAex2cheO1tRd1oNZhk+9NGodgsoEX2PzyAsIH8cFxRY3xRf
LQTIU9UJGj+bQPHyd3b9uToR6LuLOBA9suzQevwTHNr5qJBollaZ85p6gLEU2Ho8ezdUcS3FsDRH
xk/AJ/P9VNj+xI5HxDvcaF8jac7tUfD8LjTt9EuY6wOJ1++8xuY2UF6jM0LIkIrH5wcaYsJMrSFX
M8qxk8T6LXocb6jYMVYTUUrglBGORpZh7Dl+fX3FFcj0qDcftmHR1ftvD8+oyIYjR+WMX1yn8Rrf
Nb//0bHQHxZ6YUDAwVpWUOlGDyWtkVQt1Vl4mGFK56u+SkDSWZBganbQmlA+To/gId0yyK+lVkaR
oYbj8uP7/oIywgoWQaNIzH2rwrZ7+V/Afuhlfh8uidVLMCuBZ2J6G0L8+EYAffJUty4tbLcJse/O
+xYF23IinrDMZ7nEMkiiDyeu7MGjPT4EkAh033fLIJUuquEv45xc/V8d0Lr9payrkZwdxcK2bndU
3f2VnAzNlRzBdTY17xne7KIhPz5HtaYSD8vfezawdyUyHqv0vTImATadbPvaBopaaw3RtQeJpMWu
cDcAx2HZFvCT4lPv6HAktkrZMEFIbSyDP0B5XD2nswz4LmlHKT6+L1MsMek+y+JzMZ9mQh4I7edG
FQYV9sfh6t3Ksx/4N1jcv2JNfMQCT/2sbybizGaxCQuksUpnrK2kpXbmkLrX/j3ok/u/Lu9HiA02
Urq+bTdf0rkR2dzt5s7tprNLfJuoDch3uVbYRGLtDK+RQPXXPRRaK3bohZpiSP/D7TMh4sgJv37c
BaD2gCfjuwxjrwcAlg5W8S6Zpn63sQhWt5pA5aASwsrdQy8iVp3L7pZ/OiCPzimMnT5K2zwslfBr
mwpWbhuEBhnb/15Ks9Q+QT9UWdfHnoo/NBT2wuBENoilcYqFgRt4YUvxAJKw66am69Tq2VwFFtnn
bu4iCWpHiNPq2azIQYgiyGwKk14oDooXbhdKs7gfQmtGJJOIZLaab3rvI1h6T06sdvzNaAc7Yc7o
htR343rJkEPsafd62kDeEgpd2SkHfuhlMtmTYF3AYPHoa9m11WNUVkNH2fU2DryN7OTAkSZ+V/QG
Gz3IBR8h5nrISbx+btVcAHakTuCkhAax9Dz4JhhR4JLYMsa1osSgd1uIxHrw6+txvAv+5PO2Nbsm
c04a8h3L10oOK2YeFeLguK5Xt6wOQfdqfa+//QUnAMq/oyYg0iprZRgx3Wvj6wnfJJrNovTHijbW
b4U/g+4cDLdl1oPwhsO2+Na+5E6NAoF6ggjLyVCbFDSmkuAOuuXY7fdkq7NAm8WxgL3pespNL/5d
GPPzSEFniRkbGXsWgYwt+E3qABunTA6+vfih7iyhUeglIKJlfnl41rqbQyJCdWEBIHb91PfGUCt/
NvxRkK668iq8TM8OGXhqgwmh/5vCxv+H8jCLKOWJE5O7506Wkqbm9+0Sf+Us4BlGjyPrFhp8RhHr
GTp6oXe9T9bUVSbc0pRk+/I+07GmernO1IoLACtIG1eQ4XqRglJzwxxJbSTCzFjub3LcAXTdRurH
DgOKFd59jb8DvxEBIhkS8x0MotkZ7dggTBTqJ2DjXuUaUF2kC880WtJZNP++Ba38q91JvV7Y7A5Q
aJXTs8dPpBkuG/X7X/kHiUZGXPW/ZCMPZEbcSNTAMr9uqYTf+QHaYf6KDaauREU9JVZKKN1Li64A
CMdQHeKUEO15kBUP0WGQwYUWvzvFYV5uI095CuKOhhqLTJwbHz+ishIi5wgRcWz8RPMdPCRpkn02
MrosbM+6m+sLsTDcoxDRC0Az1J2fq6MgGQhYczFec/H3C5S2WOqbi1xG2B4r13HUiCpNjWd69kPn
jhdY6KBf6zyXcy4+pcZVjPrOhmSHCuz2OkMtA7h7t86KyHyIiTXKSOWSaQong+U0QTMjOFe6z8D1
rN+5yYLQRMWR7t3HxmFK+ftqJTlRfpgnX/5S5zolSKufmYEBy3q2mHdTSYB5rUOS5Ha2RLuF+VeJ
DWLIkkHKS7zRqYvkZGzFJ46Y9ZiWDlOk0xhyfC3mdGbFB+ioJAdwgnwnoa9/man55xcp7UfnK9y0
VtY0JBzayK3m6aF/VM7y420Oz57ZOBCP5VkrgO4ZIriIH7hoIeRUqXHmtGgPvODVyBGUN//wMmHR
MfEZWRCbpaGp/mZS47qUFYtNC5hy/ihGyVJ5J1kXFBvSHCaiOZaOYGKHZcLcckiDeHsXBdm0OjJv
349IKvCEastbqGceKklzOVSuk4Oc5gLeatmHx5SQTMAwXuAJ7iRrdwWaez9cA6LBx/D6YolnlJzL
iE12Cj/AkLC658NgCT0JhI3sZNhmv3KbCGPl35Cqtuk39dEzxUf9pBGZhyS8ka+nSeZw5REl+hSH
QU5S7Jk+/amlp2mveljp1RH1p6mzx0iRuK70IBolmy/sVicXkB2XPj3/yr1w3K/Z4JJDXxDzyCZF
TUk1KsBs4lD5ggjT6A8UVohrUgAWr9UpIwyP4qWHf1iSWM2Hzi3rsIhcAPzz0Hq66+NyoKPWKozK
4yrh3P5Rgr6uxCNoMi3VLnPvVEG4khwmn6EDX166qyllVgBN1AveAwccqQCLfVuCbE7JnVj8com0
71Q/shqcEMzQHWJZMsUUjkoyYj5FjnwgaLT8ZvxRzQI/6FRNJ04d8m5ZRxkL62XERe23gwSrQ1jb
YVrMlnyIlleHOoq7VzA/L0DJKl86ThcsmLuvK4VDm0kp0gNfJWNUtPL8MMaJAUtledXEVwIEzvQN
Ohxvj+RPX4jwqQs9y8Jb/f/GU17B0rs1g59lpRoLvOXhIiFnDpwGsBPmsT6H7uhcnrMAwx5V23ee
UJPrFtMPzAUznL9feXVOIHHYcm9z99k3pgQpJxIOWa7AwMwhxXvEwajFzCbn+o6iWC51Al0ghR7W
XWbehH1YYfWWemHVKYLt68+y6uPFi/9QGzXpxDLlJNFRWdhUecm9zbpwN4R9UsTkUu1AVbNqT3NF
es1weYW+PSN1JgYeOzplAFQGOXegUVAx7JOhL17SZATbieUdXLIP7BMETo+j5XajLmGFgJ67SoLI
IqTRdLluMS/BuexEiCCda0AQsMHzbDNPrQq2ZdH3VyLatMpFvHh2NOuB/J3+TR8HPtECyvL9ySAG
oOEZu25k/2FSqd0SBKaZ3ZAh53ppQIhJWCaqLHx2g6B7ODj1XZtzN6SgusInyKIRx92qXly9Zzrt
TrKt9wv13Y+wJOSTzNDlz1Z8kHGokppyIj0SVTtCLmfjUUob9sIzfUTq7mbTfxSzLT/Lwg9h4Fpm
kJiVWS0DC/D8PHfjvbG5h2OUcwcqzE/8VTwvghd8w0LUIEd3imSQL1uKOiWC0SMRgDSLO+UrY76U
dUiXAk2k25Xki9BZ5BZMH2VZO05eRH08NNuJvBHigrYhR25cdH/aSrwkmmJDH+rcRtZ/EW0oPqVz
YAgZAcOZAYuppma+dJ6tj2nVL/Uzk+JH33/ChjrE63T4+KTD6bzml/iWcHBta8rsCAxHsgJvYm1T
HKXOBZIVuodacXbMIldtw/DV8qyVvsUcrnlonSeGQkOXmMMs0PzcdfdoI+p1YpYWfLi5oIgnWO1Z
sR68WTvXCyAtY5OuW4emVqmrkqEDmVrVpJuANx200R1lRWBRyNXnj3nnRb57Mx/y+tMglJ3wCpsp
jjPuGyMbZR57Sh0rOxpF0mfuToCKMTLKNQxj2NYk/YePTqaY76lwt5YHw+MmMwgtIjRcFFwwHNRv
e9c/P5rSNZrKGirxpBh3p5ROTi0oMkyNHcCvMgBVECUEu5C5avtajRy+QTIxJ/DshAV/RQ5KNjwH
godBflAdqRk8wj6IrzwtBvGOOh9sq/ZeOtlP692/Ex+8t4ji5M0AdC1RDRrWQQ05uIkGTD9bDNg/
gl7d+UpFv4TSgDiSWNk1nWcjNjqUQ6cgSynohPc3bCZbBjZbZJMkvL0rpWdR7RCv5XorYxE2PPsk
ajlyRQnWxWGWB8YOLrOH6LHhSInsD3sPxIUk3rqQL/FwQAFnMAx1+5adjOBavOQt8grrZwCGmXwh
fHkNSVcim7PwZ5hkEQdjOvCCsAEEKobWXPPjK5f1zxoJn6QMe+r1mP9w/PUHFJJA0/cYHe3VBAoA
1wlUzFoRyf6J/CTbozduZnEjpQIWe7+gU0WQcBQaaNM3/C6Lx2gOB5yUDcPa2PBSZT6BQf0506PT
5ExrDcCrqh6G7je1OPLqq+WmD+aSeHb0XvQwJFt2HeWHgxsh8PLT5yarMzOiB5QjA88h4lACq+yN
/NnQWC1Im9HfxxtbYQ/aCuyy4GtLVZnY9LuwVkEhM7pfS2WTR5WaqzNc73Dl33k3eP9w1W1KsZhx
2z1ANO9/bfLRKc/w8szP45QBb7VDTvxdkKxaUTRkBlaQoi/G1LBDWyRH2lL/k32lH1LD9oN6G84K
75XHWnKXGKP+Wwlf+ZGEDoYD9KWss+n4ssJXKOwCCkoBZ1QcOp2ZIWN0NXsz8nkSKJg33p4HA4cO
XGdiGQSwLrYIaYdEAnzoaX6TpDyyyHXmedmDRn3r/ISC+5rSBIQV9GWI0dall8bWw+FY8N/2lqe1
PlkJWK67LESvJbxFGdpABM4Zxxoi2FIw5IJqnKLerGcX+BlDVO/kqxMFhbVvJNzvd2mOIOcmnxAc
ZOpRrs+pjzKH3bUWuAziUaFRJz8JOSneNjs7QTQe4GYIsARBdyUP+iqbvr9OrZnngHsqjmloXo0F
49UdvcS2Uo1PZQovO+hEzxdQeP5asjOcWGRZVRFOSWg6fMNacxMz9kh9zdiiYnl9u+8FJrwFuY0u
+aLYOOq+Z7hzyZaEqrmmXLv7axZGaMe/+PEC6mkGsbnLz6LSd30iQUDM8Dx9Kl03Prbx2NQylgiR
PhHSJFPMkj1N/EEJn1oT+j/dQZskyx2yJy8PbUHqpgUbT2gMDXy8ZQQVeTgwqI22QeeOVAm6H/P2
5WiCARZQtCgfOgoDnqG3y9e3QA5MQT6gIzI5UuCcmJDjUzk+BzpRDjVBFLfFddiUa6t7RihIZsGr
52r1Ou0Lzn84i552Xi0SAuJ7+BVnsXLg7KE9D3xIApO/8Y/YlqLV/YjGtEjus86T6w8pNvTjb338
i5QkYvy8vycEZU2LEl3iD2t/avjZvUd24DS94MbD+3Vme2LDGS/LoyU3t49htKcyhEjNHJVKvcEX
DJon9wvS+ppEPrq3PDy35kq2dRMzWpaOuQiGWgdYbBuGWNCpAbTpopWobsQo1qvgvitqh4K7HF8z
zcaUjuJlpHwVn/gA2HHxoFSk8vBpJRBM+TCyYIVzQ43G38MaK4xpEd1BLb3tFdqzBM2i8WdeaT24
i28cwLC6Agm3nzpThdEMcl2xatKWwnfGJ/YpaOyELuAxm+Tucmo+kT5pmaJD7hw97i8xkBMbMH2s
TS+A8IXiWQUVBLzSSg34vFhJ8HcZw+ikcMjj4rpUqxUBuSCUCnl2jVPwM79jW3u0Xz+3H+y75JaE
vyKf51trmtXhJDgJ7E/425qelg3iIKK1Lp0sNN+wvSq5AFIwgKeWC6/c+N0M4mSszSNDKjX9hDE7
xNlZ5+5wQW8jstf7XVeZjBrFIpxYdubcQWfDNnFPxRLIWigSQLdZV4ItlMYpZXSVFwvQoMwwj2k8
RCk6FX+xHg+sYQgyotz6Pi/uw4mhCyTsxs1KoaA6r7KK10mW9MDzSl3dFvAmzZewwPNl6bMFtmD2
ruKxtV+h4yOBMC4U/VLRVdV0+80C/xvDCmudLDph65arFXlnf3QpehpzWOLReCEHgqUCpn7FeUyF
XLveufkEK9N8o8uCVaAL/zwxE1FfvejsPpUBZLlm/dwUIhQtlFhIcJqc64P/djpPWkacd7dBYIjP
5gUsc5VyYtYBCV+DV3T13LV7S0muN5YH06ckdlzMmNJqi+zZTM0N7jMeqMUii/bCC3R9XwP7gdPU
D9j7hWHoq1ECPs7qyty9ySYVKiG6bB3BijHtH9jFZGzozdHG+Bfbr01DizcYO+t2/Ik6x7TXRZMg
05KQKhov1WgD0VVhtsFAVzrFjCz1SMWn5l3LS6qCE4j0V5c7Pi7tSVZa1NQv0KF4ceCSfQAiE9tf
f0LDQ3ZRTpX0sr16nFOHZteOYiTbZnHnEHuV7YmK6E5mLwRnQxPZRBdUfBxEAaFrSrd/n+10izLH
mt4NNjnxnYEgzyFkrUoNeC2otCXETqRnyQ0FDO2e8GpaniQGpZP/AQ/natXqMx/lBP2H/cghNwFx
pzQlqi6La0Hn590fF4bcQhK/P1HsdDQFjReu4U4YemmaeGb/yOGvFGgZkSxZaJ6dUMRziOHMg+Vv
LdfOrn7YCxCDAqTOp2V7wUCQGGcSfRCRRXklfiJy2UlufSl+fGMwSpb/JPh9ycwSHADGeqkPH/k2
EfbjBbXYeHXkxUXdCahbBnrAv1Z/Qr7o1F1K8P8U/Q2zrY5ITehY1xoEjNli7kXQugf/mwnoB8nx
qjPaVwKH7E8DSmqFWjuXsptleQ0sGp/sQYkc9ia1DU9xwDCQTsqewKQeewstb7ePVaelOm1dJuJ7
fCwvIYWjtLmOZFM6jhnnskLn8UIC/deFv8G5C+GSjwxSk90DYujSkYBCl1eecfOX5KaWuaoxSEna
nFgbEWVAjmpRWj68w5k7K05bur446yZ7GrDW2k0RDYOxz/7XVwatorT0Kxt6EaZ7xdWl/bKOjdvr
K3IOKjwQjS8c8c9KtaxbBBxgiNDWYVpxNaLM2qswv/CrGcnzWIGlA7QB6YOJWJPdH055myMH7/TF
uaOnAkw9sEgvUu7HueF2XsNwlDH0J8j4wT8hxhN/rQeOlzyVz1JVYoe/KON1i41Bufoi+CxaKs+s
E5914CIE2+175L09deJngaEo/UbhNd70XjNwp6GzFwdyYqj0c53qIlO2cUkf+E7dEFblEd3qlOVj
gCVYFcBFV7qp4fRlDro7jnYnwcDllD0fYi+VDSBb8lC0KDETQlTygxPQZSc4pjKhw0mA9m5eorGc
KADS5y4EBCMFQEhmuWSM3F9kLaehYisFzy94Fq9pAeEtH0oLyHAB4kdYmcuzCaw/BJN/8/2ntf7E
gi5iHkB8XgjlUVnMSkZn8mfXYg+yEbm36GJyTyrcDV1hd7FwPFMflqBTHokkohUiBgYLcS8hcL8g
0VIUJmzPjfqbXA1WJaaU8lUlOCFmBUJQZ2oA2ERaofnXOZsstRBgQGBdATIAEod4a5rDYfY2hIcB
0kvTdr+jl7kn2xG2FjQ5ck4VWsw+efxeSnW0wQ7/sED2EuWrK5U7+be5TZGI7/MbjHGic1SJxmBA
FdUlia3lNS8kKgFli6E1f7rdEhxl7Hn6hbA5baXG1Mpoz/zfCFR+dwydQNSngHBfyqn7MumUASoQ
WjxUT7SPGWgdA+VYPUyXxnXvpDny4rEdvIO3kuXAQ/rf7cVAiRAl1gmpoFD4d+Z2sezsLNYKpXUE
A8PtC1jRBhM4JKPSU16W7RSrb1+8tR+TQGAS6YlvhNJXh2RL0g0NRBUrRb2ifoxs6ePYc/InqZH8
a75p/u4YFUIu0W1v0BIhAu5/XS5k1A8TnTT3Dw3fe90ecawP4MwtsCAF/vU+dsVESzQoR3ccVRF2
Aqdg/fslw8CpiMS8mNTYuecP4+1GsJ990R7nYmylmeOvgeb0NFQyIsdjldEAGooPewKBwibQO4Ge
BmXalsPMhZ/Ej6rqtr2zPEGDhU3qwEdyQGT0KwDEuWh8ZL4IDKkakGTnI7S/fFnlVHba9pOncvET
cMs933OrkOdW7dy3tjbEb0uqeqlux5qmp1RR7MwZ3iN7VPl4j80q1EQScAlKfox+zvIPLBJzPgHt
SjL3BgEkTG5LW4AYW0TMxSZdFW9Yvq2/Os2OmHmqDtvERVDxMX8dlkRfg3D9GAZ7xLmlcVIp5yko
rq77Gp5FhLdOnxM15/KP7SCUhEAWiuEXwShSvOFzhSjGdK+R/U0B7GwDlhEGewicRNeOkSm76ctQ
4BF9y2oLpQOY5uPk5G/HzNMNLVIbF4wWguOnBeqC3Iir/biKPDSsS/II+revMzTrBI8RITbWoU2I
1Je5E3ez6UawZZ26bCP0W8lJKzAyK6jpASCjjECdTSMyXiB+QPnTk61JLYdlT+FaEY5bfe2x1Jkg
B6gcvcrsRbE/Q5gAn2EgRSJ2qqvCu2Ti8b/F0Np1Y3nDIa3Ps6wmNvIsAyFR/jf5BrMq4v3eyz4/
Pvhsa2BTaF7qhpqbAlBI+o25rouN5T4wHvkFe9GcQtZkzKd6WmvvSnuUYkToOf8U8R85w2LDgZe8
0zqZmnRoKTu50eLNFhJOl4GM3yh+yxtG221EJpN48bXqJXZ+2h+yHKHoWaMkZH1s24rp7lV06ePF
fITHTfymB7h8TL43Z8UpIE2Ae/Q3aP6ze57q22LWDqIQ34mhSf5pt9BZo/mKGUv8m7ECeo0TUXjV
CJeBLMySEdVibYm0tijIO52u92a2HCEVTaxvGvGS+MzUOxViNd7b/sFGAv2hzvLE8xACq+ZNAnfo
qE/cK0p7k0vuysCodLHt53aPet1a26e8pfAPfWhkeR3iIVl51YwzRG3OSUjsdIPAdJP/YL0tK6Aw
leQq7ZLslq8dbQooxP1KP0tBz1PBxhh2ICRIfb8fivTbKJWJPEXWWGEJfPXobeC+cn8zhcp76F4l
pr+Q+PX+Oz0+v29swuP8vhgVJIwIl0d3w7hQwipPVBg4AAxa1KsZamonDf9empVio123R4cGpj6I
+EAJ3hn6DsMDIdb/Csn5RquFDgPIDckM2ftfiFvX2lCqxp3BsLC+Um5yhKyshg8JU9XU4CsB5nUo
aB7GltWjTykRDAo+oAW+6OCSan/age77SS6hE31+8LCGdO7nKGZEwOjUN6X0Wk2GDMOHGT6VLtBp
HQyE+ogP3miBlGEUCaOS6/txDqgeb0RWUd/z/FqJ+GdUxOoEcQxD2Y5a48VOnK1gfDpCmFrkzl1W
RRGbbfttKtc+DcuNlsUWD19ieq3d2T1CnyExpPcrmDZ2Ij/WkXk4dk37b1lEov3IU4L8yHgkVTJj
6TqeBmmRCl9af2LJBT3qTrWd5oVlYMylH/t2792V0FDzbsIYKfzJNO76vUE7T8GykGow+3OIHUg1
WP0MRFe60AFO1EGb6XHNeeYfdL+m4LWTXEHP+dVI5SxrAvEvqYOmUqXhiPLZViIqqDl02dpzBcHc
5qzxNFG6M0EfFPJnrugZglTBZTCNjoOcQiIJHbX9HecxDP/n4PnJKG93nMmgxjl/MMCEB+h2YfvB
0C62bRgRVPvb77km8XedlGCOFDiWgu72Me8O69RnI/l7Rd3gXhmbGDHTSKnQtTmlHPG0Lbs+TpS4
F7Mh9X3pLngNjL7PbSYhLutpuYW4bWfmgXHWQRqrIVs8X/jYwigmziCO9X90X1QCojQ3XIWY1o0N
fFg1NmZ3mOetAz5LJ+io86IuTr/TmwrjC1D6rWP35V0h0L47quZZVYitMqITmgPqoJ4Vj7kK5Rr4
929GR63fmmR7V/T0rjc0rwThjzRSvYxjC8QqYgHg5TxIOknvOGiN9YDlFpbVigCSm+/xPlm00zUi
Adld50qu2aZmMRE+q+x91DyLkYhHCyl9SZLjYVKaSCLeRYDMmsn4uDWCUSBm+YABfh/JuQmjL5qe
5t8CPewYCrjjONY6GNaVAxDyRLpGyfQwg5OVeqOLhVzZTUfOj4RGDX1U4W6+mum3CvzJ7NDJo8m0
kidPTm7B/+3QRXwz1k3BZp2c2MK882yg0GLzd6IufHSLOWPh13ha/KhX4vivhMgoF96iPe7fzwv5
fQHbJocwQoE5B0aAiTdJ3goZLKedXVQBtoPQBxjn4T8xKDZercZ/QPIxIlAs9DvsRoMq6mWBuscx
DtPDwIo7UO+p204gVe4XIDpo9KIIop4oq2GBJld5uTbSBrlwii5fEHdWTPkARyHQEvA2g/7ze+Lc
wf9KfRqnim0f+lq5qkfWublI4DXcp4m8LJb3NfiBvEmzNa2oqR3E5mrz7GVWqJrRtsi8+KeKJWTD
bBrzHXrjjHLTfPwQ2aThWwBEY0pevWw9Z089lbyoG6f/6d3Ij/I3p/p1UhNXVSdq5kVRVWsqY9Qo
9KdD35uiAW2bcoa7E7mInizJ37+zTQZG8bE2TrMzdcr5o4Wetd/nYBUfa6JmgZQ9VgwpSXBZfKib
ETZmFC7oe1AXwnHPMlIb9h92M8aO8va0BQl3t7mWE7kitb87g1txAB6XhtdRlJExWzHiuD2PExdL
ICVJjG1K+gsGZCJ+f0DNqhTq7SEPhJw=
`protect end_protected
