`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hClBRqciFoqpiW89VTtPIYB2OW6RZkXsvfKlR8/pV0rDEJ519AehtHrizAojBqwPC66Phbah5+QY
rq5uQvbDyQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PK4cXtjRFS7EHlG7EydbmTQphhPpFjMpJ4TvKqZz1Q6qxwGUp15E4C1cQnt2dleENsAJ2FuPlwH8
0MS9idWeat0+ksi9jOM9EW+Fgoq71m4PM4GbO++fPBk7z6V+QMln9IsE9wJZyU+0Ji6w4RqDiAQn
JUYeIACnRakLrew8YGQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MbhlpKAz9aUKZP/oYGMbhjJbXps5w8sKKeFNLqdZyaOjBZHRHS7/TWkRZDVRY2DHCUhg91+oFtqQ
u6QOp9mCyYRir/u+S7P+7vX+K/cMJ/f2cb5ClydKSezQKZQanC+x3DMmeygd54IdQ1uj7UxoUbDV
II4jbuiF62/w+iBzibMQWC3wxM2Pz8fxxA5K5P4zAiEu+xGjKfe3QL+IJAdm34gOdyT84q/2QP9c
/MzZA3BcZBiIOWNOaWCqp+DRiRub5x/I9Z/H6P6/tAyxKk4PnExuVp9XYsrNbUYJb1nyGTunRnrC
S4JsH3jCHyzPaji6Pzfw7d0gIcAcRPFXxMgveQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VVMqGkMEbL2lQlJUd2ou7F8GrCJazHIoAV+Yqd1OSa/oPcKciUIJe3IBaTlI6J7TlX7b9mGyCB8r
OAbLMRADx3vvuGVCvmhykOW9jNokxe+6rIaJuwu4UJnU+mkA3UTM/wVMYyc93l7AafqvVvw17KHo
jeCNerJKvvv5JFD40kI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P5iIFIHJUebrw4WcHdY5lRu1t2m2j+Z0pxQBKLiEOO7HAPdtVJkh5RYUs00Tefmx9XmNjbFTcZmf
zwIFIz2hkwI+4OMFOZwTrEuK1cpJ/FlyaxAqi03uCG+cX0zmg98FIpHIhDEzhZRYZojwT8YnFypO
U3l/ODnxyAShz5kABlH/n7ZZ/jiZ0kLAzz+OU5+JBX8u+cVBa16Zjxrzed8y83QAJv//IZ2DMCcX
9KxhBoLofdkA0+Vtvn5kb9n7ptEkp+wZGAkJdKu20PrJgpE0F1ELCb/8XSlzrXQNfwrn1vMAnGJo
EF3e9xApiWGgvNLQPPKWptKB6NRNm0iIzd+k0Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8032)
`protect data_block
g+phTx0cCAnFlOXaESCK+g1Zn6/a4z6kVZSpxjFfGes4no6gotlTKOMOCKn6sWM5UZUlWWXhGo6Z
NUiykxrLeq1o82SPlErnUNDOFxRXq3uNIhRGReaSnz7npyqcdsf1wd5VbX8XZUgc8q/qZfQlsoBd
4J8uU5ASccZIPTQrm19QzL7PqeH4UIF0OFKKR87iVhtCgXAQFx4hE84k9Xvo7UeOf4R87CFgCtyh
V/Z76W4RYgKBli6gtue98yuFwvLvvo2nUanrXT9Aey3jbtUqyxu3lFdKxKQiMRftfLdwZOe31Iug
lTuraT6lJzN1XMI7NjHvNqAGuIE6XpL8WR00ClRSj2J9YFGkC2+MjCYg6TVLS2hc7Y2PtX8VkdU3
usoZbqhk0gb5hzffNLe9x1N5GzdSaY0kJ0fxjgA5LG5wmij10smHAHwXjPrzFzjgDF7bHtKw4O+h
/BB8kTNvSmu5/gSRXKb/RVLrDcxTmrd07eHzSJrDJFsDq41KxpW54gScqmY1/WzYoqsx7dSVpGPE
UaXCMAfU06JTxPkrm1JpVyZGzsG254OpoIzGSPAFGkOkK0+6OyZX4lsrN/k3kKOEANem1qTHeqdV
XFh6M8F/zknZseg5gIG96ry/L3K4fsGOruBE18m77Ei3txOLH8Mw4aGHF7DSialw8TwmQAVJoUa7
p8VBLCfRgptG8dGLjk4FDON6sfFHgqjebQq0VHHTROZRSHFm4mzWEM2zjpohKa44lxueLYcVVmZR
HuoZcEI/dO1Tx3OlKxPcODw5HDWgKLraItNqdLQzhlPtoCaqPSVESPxlCVqS9BfbzO8NxSrhBvlF
4ITKOjlrYbnZlBOGcbl0BjU3MoCIoJrc6vZH6j995doBvZnelxppKhxeFjQofPcw1yVmTTWLfwEK
IP4SVb5L7F5cbHvNMV/jc5K/vjJVMcRguBTrnyUM97XJUCIGRIbJN3k/LMkZklwtj9JBfaPQ0R8F
7QeXtbUW2uFB++TwQiSrImMaxE+PjFkshy0gDv4IpKYamBIhQfKrGnPPCsoXkBQ9O/IqTDzlaLfC
PC6KDZmRZkfqwMW4H8F1JuvASptcgut6qPwAtdWv6xn8VmZIfBVkBphgkRErWs9rqa/2AgtTGAPX
+h4g42eTgV89/PLJ8LB7b0YzzQRIZLmT/qtnZI/AFNj5TQau5vwsMXnC5O8RQVamuhVjr3MjaLtb
unEV6NGKET4dUWg9dcFQwM9XiLwD/oQ2R8ggEoNOlQgET6z8/81Qx6N4g+JzZmqn00iY25TSVAwu
uZbhZCdBiR32E+Z6ihrVkSh/AMIwpUMiYra/YLr1JwWzRSi7k8LITXA5cqcJd/IYfGmmGVxnuR5u
RWZLEvIfhRU15mvzFVjf2tvEm+6oygu1lbWlmZ7w3aYnu3SEipHagG2+PjTcO8V+eJE90H/ytRJF
EmTDmmgq4WOwuNDqpBnr7vx/76+oyDFlSCiYEsyrEmb3QAknFFXD2Jr/YdkBnc18kVme1rccPtt7
itaU93nKvUHBrEgXlfvR8cpT6S3sSsoigT7P14aw2AOADp3JntWCMi7K5IQhpbcjkDUsdXvazCOY
Cr0bgqVYkcOJE/wbLHkgpOLsMiOl6ponOP4je4y/V6fuh87GJhH85erHTEgMUR5KNAmbWsjiA3xs
w1SUag1J9vCUE+K7jCSFLJl7lvuKOD6dFZIXRDrlcI0xsuMPj7Ipb1Q2GcWrUM7i2OkXWAsXZXzm
R9rm7rewb24kqDuZKrUNq3SIgCxBzEGz+LCWtLRqgxA6GyDV2gIT54Cw9KZ7JirYDSvBKKzB1nsm
7mQqTMVNCGtgqFwy3TI8f1Z5yYdmZcFgTBy4Nc0cWAyefV7xX2YRIa1z88RptA7jcIdJvcgFokSe
yB2gomn7ady+iS7kxlXhsJnIBunWKIWI2qBGSE9zO2S0/didi4WQBJ3VRdNoYBbXTC0raFzOnXou
q+hFoFaKwZd801PN8lwQTb9Tj8HJPj+dhzmDxF6NLQOm4CcusWl7L7Yki1vY6uObxjOrQVppsX7k
uwau6TEAuuPGZkaUPguRqAsCXOlXdukt79eUl3ffGm95aAw8JjU9JvE7OpNjX8TEVgAOfKPJXuMN
QE3rhkE1R7UFrHmDJdl8XWjvG6cgZbRD6UrYH8WKbpRaYsmD0qOFwoic8i08ITos5HgGWE9ZOBoY
smStojIeLJlgSEXwDvtUHaerS5XRrjPs5oWmqxTkp+4aLdq4zXl6me+fF6sfnoe7P+F8KQm1vdxo
coiF9zOPGxdogC7XKpDQyxpgR1z3YoSxcC9AKW1/6qOPunnaBiMZtuFpFIBq3uWy6yzc5u+ua7ul
ekPhPR9XW8aAbDyl01qMaY1lnlgbMJmJ3LBTc8+WZRZPUGoIO3KcFEIsSH5kZUNA9P26cMayvfN5
XDPPPgV6kCNZAG5j963Kjxv18+NNtzA39qu3SDLOlpN4OsbYaZJooRKZrecBW69hRkUmaz8WLFKa
VkQZ5J7lJO/LnXOP2xvOROy1QjYcwwYi1E6lwhzk9xBbuk8v0Dj6lwFAqt6pg4k9qjDJbjI/YQOC
AqteynqE4c6oDXXMcr4MdSl42tEpz9Si/Zm5Mwim+EziRgwZzb4uoHBwCv0GhmtzIhflpORx+RRV
tUH9P8jm+cDktVYlUmK2elGZjyODnYr9z5/0J8GkJ00pxSJDWP85G9g0OPsfGC2ebUT/tsLXI/WA
xAGoeu7THrbDmoHI/6VYKUtrPVjgROvfrZutqlbqI6hma6zLBMNhvkYkzvzn2Vn7mgd/qPG/2bUt
UnAyx3nT3nj4NknLq11/64bTypbqsCnUo9mIXogEcZcfoI2eQtuEWcQv29z/nkHiQrzeFyBCid5o
csk49OzFdzAyvVPxFeBBoWhTEuhkDRTti95JLJoAciGLM/A7JsZm861j2NOzFEQwZnYvmb9tDibZ
hT8DW9BCv4nYsQv9ydv7BCkBzOnNBs9akluHqOL1ZEnWGF9c5PErk7V1Q8PS0b9sKRHzTg+IHGkx
lMzSFa5AbDchHwhI2Nzdj2z+Om5GdsnKgiFTBtdJjL95oqNiDo8bnIAAGDDdSquo+/NI6tAcGtVJ
XMgSKdOlJnw01PWmyisc2XqDO3z3bJFnmfxsjOktwvkCP1H577lCE7Am0K7sHdZsdjn2onGsEhF+
veXHPqgKR3iHcsVxrg3Eb7Gr9DtuA3MRdQRzbhKa8xrbdU9nzdJYfEEk5J1xR3jDAzJkiPo+2gZ4
UfIvS7RssrmK8DQUbxJg7BU2ADwSA1WKL1SRBerbPu9H/6aQJUaMeSPIQyd0zpZCvY3d8LGRarGY
wK3DLyAXTPd09onpuL/5HWt7ksnMDEWWBpZbG4bTNdLtowK7NSaqsTkGr+JqyHKyQADNadhaDGiL
OhQ/PxHgX5+Mf9BrJ9s6MGcXMx3Sbk+GKgmyPbobjlOVRnyeBtwkdV+CiXQL/W9tNAsbfRn5DNkA
5CHYJWvpJfwGzdZJHK4snO4m/upar6hpdOXU70huqUTFKCt8hfZUXxG7Q9v3u3WhB3Qptxm/cG8O
7FVRenXr0eRpXWTwSWeBVlI6VWCFr59dvvjdWUcMW9Bq9x44DrIQBq8P5FxsT83Kn1tzZiy19Ifg
KM14HW+jWcS3AejB70mBYDW4B3sq6S6JnjRIkudWhhSvIIg52iQvdSDSeCDWBpd3sbzm+UkKRqXw
YVLkJfx6UncM3Ysvcy/bMkmXf7rDbQebyZjWbSrkhF0wYmQumncw0v7sfjt/9pBgz+XDd3qnIZfg
AkJEUWohqUcBh4mhqzBRKNZTBf8JFwZzGW+m2Yn9qyfQOIWD9Ivy4/PwIc2oU/CBeysEGDJdkXUS
sYLMt0ZPLk1elG+Al7amFYa/++QicCBSBlDHVVSPHmC+9oiGL8Go83J+IDRNqmhruo3W/geV24K6
8lZP32Ots5qnyRrAYNdmTtZnZlI8OYvQKOKjKeA55CbN0ram2jgDR7k1cwsxkMPVZvlnPSVyyCHp
1N8nNPrp7B+Q7HjsZ7ndKPSJ7/WI0GoPpi8IJyKdbfNxp4OcVaOZvWpAuhZGOr/kQhEfUQdP/zyz
5zLpi2gh/HnEvmjd1eftDF/GelZcaSvSw+urTaUS/Lsi6iiAnefqVk8LlvQdD/JjKzxx8zsFKlZe
T0A9Ffzq/LmdtCZNPqqlKJuGL2KIkyHbCPhmniEwbh76FvrThuzdsp/FBQSM+LXvMMqWKJbDbhDw
oBnxdM3WhcB95t2rldOOMlT+fYX0zOzblET55jdOF2+6J2/4RAKfUkiAaTyR+Ivdk/0IfxvvtR8O
p6014CxCb4GLrsHoFUrIoSm7WoCTJ+wOxahMhcPNABDUOYEUYk51lJvoq/jkYBTK/l6ySz4S3j5x
OWQBPPvOj94luhoXwjk689Uzlu4ulBRtXypExr5+JUhaS0nlSgoxi4lyMC4p0A9vY2p7cxL0uMFd
JF4e65DAvRZs4GNvkkyXIDgkWOkV61k0alotXp1KDKVkiQJ3B6PE4gjjn+H7JnwNNwnq1NuOto0G
rbb8lJQbHqqiNQRJpiH0k1+ABpdXh2rhYE9lJbJvHM+BWENSIEexyQg9MBAgYmzHfuKb6njOP+8W
Ge0TYw+Bbth/wp56D/nfj3+PTdsJ8wOOP49j24z1Bt0a4yWLdG4vqS+Y51QHwUJfj5neYMzYLsf0
b6rnXDNdWh4Prz6Alvu6d5L8w98eJVthkb7KSwnMMRarn+tkslPQnwWx02FR4Jl7aYGiUwMwbWMF
Uh3Bp85IwQB1KSRa/ZiWiKmGZ44gbBPwRF2caUoF+qiYhDZe0ZEOs/E4cOFCBEJ1+UlA4XAOeMWK
S9B2FZiZYiO2ufkr4oo2VIewuT1kk/Xh4w+DNUZrpocehEVbFjrfcWF0cHh5spLdST91f8vxNLyx
Rrx/J1Xgb9zX5DB+QbXfm6/A0+8rDPlznLuWxaZis4pmSwI1EUNKMfKmC7iZF+UioaW4YZpCzyn5
nu0Q2yhOxO7mWORazRngrTU86J7InFRGGKWkVOg/LhSC4p8YncFPX9Dw9ABiHBrifejOKDLO6KGZ
AXUB/FD/Au20e/1d6TKGKnVZz5PnYQ0e0SKYDc8zbxR0hrrCuUEEi/Y7IPuklGchvzo0Ul987Ovp
GIoaEbbs1S/IMTjDQaoNJRaTOb6sS6h1wCCZ+g/lEhh/YQY886KQ9isu3/7XSxxM7ln11I/QaDEn
0Jn7ElzuEOdgXapX4YP0hrDFDIgmFX5xbbY/sG9dJqQJEujWesU/4TYaCpmOD9eFhKbRCnbMXN9f
bmB693oG+dkquge6fTeRsgdSUSNXo51n/5Kzr9q3hdzT/UDb81j1grmwqpoCSmVnWjdFdviZNy3f
HVKfWXHRZr6PD1gJBghPqlO75UYsTLjRIGCQDJLcNUsV0Pjr+N1Tk4jNlJ3xcAIW6g04mKHMRgfE
J5Hx49TVF0N/yeLgKYH5QJz7FEyhSznMXV5ZU38kj313cIywbEFlvdswJOEa43Y1MI+T5DdENPsM
cx7FrKmsQ6O+Dbx8xnMM8ftEJq2DwtYK8Ajh3MXwjiije+0ZfxLk5OMiP6xpU9VxCWe0ecazgmWT
8mvBXQ6D9kmz0Uo13tfgzYHW5Lia3eOq0epwqYVae0qRWE8dUsPmNoQr0Ufn+s877aNa1zj4928t
Ilw++If11X7+IkaR6KQ12vZ5NbHFl/IPcMnVRtvGk9+dF89XAaTr4neSWhJS6qZlkMM59qXfz9CO
dns3zufdyPtA2V6WyrloObhTk1Sfo8nU6lolXZDCLSFKlC/1CMZFbQI6nKechZ4FAHxH5Bh/aG+o
/oRTKAiK2BYdfjjTH4zdKFCgg9Ql7frD3D4nKH1aikECHD/2L+sAFvm4I6H2bj1khMQuEJO3jcmu
Ikg3xMbOop15OmA6QaHkhP2/bjp7GGBVxt7+pDF3MFrFzw0bbK7mgyizRfCop7qRtnEte0wn0si7
RJ9zXzz9J5mMoIO4fk8ZrxIE8QBt8Aq808Dyd0QZ5fb3jZhrZJ/0NZAvIqd1Nysq/pP2i0eO7mdo
VgCHCxBtMq9EBJcEiR4zRHQ+jp7k06nen6aw8fRImMRJ+2BhhCjzStvRhdnyPGKxsvj+VM62gA/1
oNbGQq/zc92hyd1SuCIBMKHDYIYJekebF0bbDEyTPbIYWWjkFlnKXwxTBlfgRyBzZgDdYzbFqqlY
i/ZbPQRNZheKFla4lwN0EC2z43vUiUnSg9OMIRM2dYC821YkdRgGZCi1/zYkkdBMImLI9ikFsqvF
fHoCzTphwDfn717qypg9ZBqGQkKHlob5tia451GLjGL9c587w5DxEDo6QbdaL4lzD8QxhlIfU151
Ye044FXgk/yGk3DZxA/IB+FmfRUmmao0i+I+GE5XjH4nk7vLMr4EFl4HyI7s0mZErkMjIPbTLsi4
flCOQdqW0mdMbouC6LRuRAbiEvwc/uBjBPLFn9+kK0jpzWJD9s1yG+a9OLmUro5X6EyhMcd/ObDa
CoGzl8SoowY4jJrp6ZCNypTYKpVmc4JUzcqluNMz7rg8UsAUyXKIl8ztSkoY0bQs9YEgquxFVOEo
s4pGVBk+rTz1/SGtgIA/y4QpYXIcwuL+f9rObRNzxbuZEo9Lqk4TTRCQmyX41eKjaeyA1kmS7tVu
W9ekNmC39L7Rx853fWEUwb/ZCzwklGBrlAuyQc8nysbCc5+cSNYifGs0bx3HqAW0IUCClbLai10x
wewQy6YRep8aFWuKAAsIcu0Q5+77hpBeUzvnWo0cQEesHa0lmnnn4SwRKXtoJ5Yx2GFytVD8Fbwo
okZ7OPeqmZ0LiRh/Nz7Zboedi0wLydHSTPI8RIm/JZpo2xWh9L4kbII9y0qczBUVapmzgyee0/UE
XIQoVAVveAVZTH3YndsIRG/EW9PiGw8Va99Q16biC4oAv6HvT0HEA1NdhWdwKpc7Da9jqAI2D4Jd
x1u7MvCw4AhUeHdfmGMpcfd2UUqpFfCZ1pHyvZxjIukXjdVahAp0+9hpVph5TYuqmZa/cfCZZM/0
2NFDameie1AOT1PqSOrul9KadidZt/aRGixS8tb9UIQ7qICDDvQzLgB8NXHR8Gvf/8MaGpuevTAk
fqDU5WqyONN0uFUVarKs9b+DSz5HNDtfHVf6w6wEFQM9YfUdqLklC5iTTmzr9SbdGyck2SpyjEQg
P6Sd8GF491gIZukbGqljU8p/91CL3PpM7Jp3dgj8k3cNnPfJQNA3IQl6pSULCTT8Jsi36Ni1e6qM
+VuhFm/8Mzhirr35Q0liNCvYcaJube43SIDJ58xCR1Hn5ZX5Nsh/Q4Tn/KUV3d1l1A1gkd3HN48j
fJDZxcOY+lmcsNt1DO+TeVgvboeTxEKDuH2VC6G9swRzdSAVkFAeg/z2/rYqu4yBwubRthXL+64B
EsuKMugcZIP5TQBnJ3iCJSVeojk+1QigCt/Y/MmSJ8jXlr7jtfTl44E7kN5BhAPcPhYg4xWPelNO
G13Lg/zrBFOAR8examJ7QdDmWrdr2UIJyBDuniKPRVI+OMpUf40M9QLVSKF7z175MTZca4v4ZsX2
dBseUQ8ZzvlHnvDGBTn0YHoFE0pKQ0pRk9wZdDmlYQxX42ZW+WCKbnn7CNF03cGiM+dYNkE0SRT5
zQKdNdzw7YJK3jZNeBy9vFRG18J0ug59TrbYq3CpAeZdFC9Z5tLMBbZeCXW6m/muQaevxAXbLuWu
Xc3ocdvEFZ4wAKwstsZae1dus3wq2s4RNzDNQThdtn6AaokeeDOV2HBpMfDv6onP4ZNAQ9m2D5Ht
BW/BreE2/0LYNViaz17j97xKShujXsGX9gU4GVNbazc4PE3rBXSMb8+5M9NDdCjMTblsMfv53oN8
+BVEvNTpg9avaDkZhkK91IFPOSp311BspzT0xnB5+28hZKlTZ9ZFmlrBMhDq7YCAuSazNLtMRf59
+FoAFg8bSY+v++gsFpWsohky1zggCFNhpogWzi8RRtk5xDVvzPhWCZc1yAm+svL3DryBQQm/muOP
yawMIAEewCLwjJyhMikTNCBBcWCCw7CY/+zImTCMCnuHMgkIU4VRk0pNqbyzChy1k+JzibV0HqR/
oFg36tMHgDZTDVHSFJF1P7M76+cpYAKXuZ4GSkEcpwe7g3dktWWwNnEF/KVq+iLUf6y29FNdrNXE
+yB5q0BuDewKq8D+paluxHDSSKLdHL4Jr0N4CiwbutqGIIMNXNUuFF1Jr2DXjrkbDFaWA0M6hLKc
goRqNIj7+QxUKMk4FOxZBYa+n6r4+uDOSPZ56AMdMZCgBv0TIAxc/g37lSSFlCofNDPlh4BnwbqF
47Nz2BqJolq57A+kE10+PgdqLlOdH9i2FZ/5wr60VlbZsVKXZ0s/fTcAwGiYMcDgUnDzyy8t3Qxf
w80O7rbcRKTQXfZDtqYJO+PhsufM7aQB4zlMYQGhJNjSlDJbC046Kg54VDtaUuGq8q82C7M3C6Vo
3Q4mKv9IX+UztI7Asw6ABMEuO2GMP9lt24a5ezJhWW1Uj+M3ua8UVaI139Zdo7WQCrd7ZbBQULky
TrqmDCx2ylT7hCmzjMXEgxZUutP+o7bZ5AMnBqcjSuS0FABRsqZz6ldsoZ4g3kQiyxpKrn0TRwnC
Uthij3xcmuhZQMhmcbZBrs1UX6+rKVYAishFjTjCW06dPA7k0x1uigZKX1ff50iN4X4qIxmjjZ62
E1qkG4M2sRI8M6DXDWR2DYzit4IgauGXLTnSzvKGBXAb8dso5VuwAZigFMV/PT5Oa8nKkxdhqcBP
aw4rlm76WqDigcu9C0SF0qipNEl8zvxvNgZyyHe9s30EFWFayQuoEs8XmYgInUVjXPiM1+QqmZvb
Tl5W/rYIN5qssOrp0Fnpd7SLPUz5nMC0Lvwsk/7tN5t82ESlqc/jyoJ9YHehyGGD3KmColpP6Kor
3CycrE7+CZGJZ5Hz7OPPSDdBe/gmQhcKTiWH1yIHRweqWz76jElAcXTKTA7qdWEyMsZ112bxEM77
kcbz4/ghzaw0OT7Usu9ErKQq9P+JmmYXq20jphGBaV23vTFv4+ZV1QpPbX3TPEttNl2B2ksYJCA/
Q9K+HfG9aBWEt/ouBBCxZBsVTDqErFWGIzOeC/zRP5CSuD5zQvPxMAc1vsUIIEXHwci1H3iMO1WL
CBiPIudHniBDDcJ2SkwkbVF/a5/tjIJdTTm+3+yazrWAT+Z2bm3v5aeBOG3hcCODDX1O/YvutOxc
9pfmyh7z47qjJqawTIQfi99nwdhibGAeU0BD2VtZv1TjANE7Tl48kfh0eth0r/781L/voeYTuuWF
tfd6CC8IJoPVVrZymUYhX0voVvZB21olUvnqJraV+SVNj1AnKEKhP8GNJvubhqL4mjNOg+AIH60m
c9PdVjWg2JE/3w5k+0wFRjMiEb5SSD/eXh/uZc9JWKe47WldKNjKdigHOStPAX8E07k0Msrt6JX+
qK4SXNtbkwpFA5r+PdLKgjypedza9Cir4ceAEKOPq+F/oAlb2BT6SQ/XrdGDh7wo44xXP6AisDZa
tIMpfHtSxeyvodS3+oTbOnPZI3+XXeAMktZjcA3s01w2Sax0GFUvMJ6OSN9JFnvYHdxyIMMfcdJf
hB8kg8d+I9Q4NHdLf6v7sHa0ufSOQgRsYyU8WJFZwcQe4Dg3MGMcAqPQbW+2MDFKNN59/YHknIPw
G0aM0OTwFvM3rHXDiEQrUuxWIj/zj6/s9maa+1ctwyf9v4Kq2suyZRybCC/cEVCCH21poKVuG4wG
7Ua4QBvd2of++ICaXVTsOIUcafyiRmwbUSR7KZ9WFKtty0C1ueZJQCprqJkq+ItOpZzku3WMTzDX
E9t1HZveNrtomav0h2jAgz9paXe1cYsi7WZgfSp5dEYs+1kYVylpdPZfj7jHep9YC7G3PmuL/3Ym
WM8FJ2XD1+KblD5n3yz2uMWisSeCBciDErGozet8BYwx89uo3E/DVlynmk6xLW+4uk/h7roRRkx+
no7WpOMVKLW6/SZi5w0yy9I18OdrVaHlAWieWF0BN4+5D1Ee3eb+ojOLzfaa+FXuPTiAduYD3DhU
/1PsEIf/OAu302hgG8U3hWY/8JguM1TRbOaos3r6yiYODNfF/ePD/VQgOcup+oSvKaQV8vUkTeRV
Xe7dY94NC2Qmcy5lWaU3J5DxTQTTecWVgjVGdUmG4f/Y5XjBaXiB9ledk85G7n8Q4q3aU10OfKgK
h/95AP2jbr4Z03T3EW6uHDA89ASgz0a09uJXPzfITFyVPUyldaDxNIvbeIdyVz9VJ4RW1q175fCJ
9K/a6IAV3aAy4QF91ePswybBSM18U24qJ1K3fki4R8Uwqh0a1hrX1QzxigkJeilaaRhnSdP8U4nl
GgLmlSeFbHafS+J2le0fLhUuikEC7BCG+Y0IkHmpCs5hD9Nhe0nuGa0C9AuLFl/AWsUK4sFP2+Cp
RNVy1RkjtuZSjLVDL7DYLCuDQekz4Kpx6qC2QPRKv9PJkSaCTkeliOEUwX0tc+sSXgYzg3beE7cm
Duv4GCowSC+aRW8egDuKccQFcon79Isqg0QyWloPgVGlzHWRg83R/0KMon++xqq1YbJRSvBpIhhF
V8IVzmSGJ7FAoaB1qJSFkPySDY7hcpsABJVXosfpJw0v/n1zWyFSCJ2Rus0Zla+10DyEEw==
`protect end_protected
