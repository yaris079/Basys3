`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FLBUKspShcCna6XEzxM/98olEUQyUUS75nUUqJGNCqltaz2y4E+ZpwFqR8ay8BbioiktbZW4aDkj
ZbEnXwA+eA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FQBuHt3D5bFHDHZQbrr6C3o5d3G3RqURpkiYlGN0vQP5z6XFaMXIgazlNZkH5dllhi+1r/LWKcNd
/U835uYa1N9PjHZgEN2L8m0YKEOVbbbi6dPaSy0WnkE/jYb9X/5SDvVAFYXeMCDeOK01fPU/0vf1
hjupuoMeAUrtwaJHxRA=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
q0+5QfLz0kYdI8xaxkg+KnBSfStZkeeyPko5+fSEtBvpc3zYnszEJQepNIi23UIMTpea1lT7d3qe
0xadCbqF2jlKVRR6uqwdvcIGfp6vhMgNiSq8JsaYBN4oal1U2I/6VYNsOmH8ptaQ9BwqyhdAWd5W
z96rBGqUWUPGdMMm0s8TyhSU6f/HLUEA+1IDf3DleKue6TEZ60IRbURhjsuP0SK6vMzVZlKLxy09
q9RLlJM3ETWvAMvFloSmiRkqbR0+W6cuC86QRO07Aq0XGnxH0f3r2GREf+I5k71Z1mHiiawtX0lJ
BO6TOVRIdzdD/pUA86oMLv+gLmoF4e1ShDxi3g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4l/r3vfhUQu5o0WN2i6ZrpVsXdIgqo3llK1LywImsTUIJ7bGPfe3iX8aPlphPFOB4diIZdgek+7h
4NtlX0H5+lBESv3tiOBFf7jhruhGUlwjMyeyo4atc0cC+WluLoevSopjyFnBqsj1/PN4CgrF19vb
D1w/4tmwAx9Bc78VoVk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fSspNN8rgNMaRzAEGuin3op0/Mp85ruMX/sEl5atYT6pLGZxiPvU+ZB7+28Ii93XLooXNGRSK4Cb
D8FwkDPZLPEzFBHfl9E2XmgxMaIDXPUz6o9O1G19gD3T23LXp0j0ppaeC9Npi1T6Zk6qgTCu/kjD
hLWpWtgAw7SkcP6W2ErnX/k10UTurTiPS5ZGVJdXzAQLSx4U8IkdTWT12QmI6GuUBn73C4kESnfm
WQybk26xCQgpbPSnu7AlJw4XXoa3C4VzqDTSHaPt/8G/R4k1sjIEmMTR6+d4YeyZPi8rsOJ+R6Sr
4jh+ppRrYILbO2vxnTkJf9JpKYPwvsUaKKoMeg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8656)
`protect data_block
/HtKO1Ec/UJMKpUqFT2jMbXpc1+qNwWKoSdoud0psJbvxtWhLInu+RnwBztbClm1u79fW0uLYxOV
YkKSkJScgZsQIw2BvY5x+gR2JUgyfOsEbcOpJHB9Z6ABczaF69y4QsuY7qyiHxnk6BBCOtpj9vWH
W45AzRC34p/dqpuvnjWZAxQVGXL7At++An5hg/tIikFV1ucCvkTij9HGunD9LRvPgKW26wp4x41n
mMOPwP9QWt2i3xFlb9vwfBD2AllULicESCYTKlAkNbW1AsfkGOdsVjvYArLK1AY8dg+EZRJlqow0
QFMUCKJ9rZc72znyOe1A4Bv1MhczQ9dFdbbRWOerzIvdlwEXqrwiZrdj85TBdhnm/CeMovuPy4mL
mXxjsliJ6xJ/wQVnwmmvsp/JxvDug4g8eqzWR27vdxni6R2zc4FMT7CpXLi2xKjBwZ8/7YYVtnjU
9pGR/C33vNoLgltPYON25sldtyWbgRy0H5TX/a4+vE6TDvKBme4WVNfdu6JPZWQEfPhiLpkXV62u
QctbkgBpLgfVUWMiXKZLHKsQD5fWbf1Q00W6QRzcPhjnn0k//9ii6QdPiu8vhTcapOUYdPC99i8t
0R6McRMO62kMesvCpz2j02tDAFuaOv31blxjWYMW+MmKLchK03dGbzGMSLG/sRlK2akeMkBIlSG6
vsHPe7j07O9Sy9wro7gNU+f4oqO1AQ0yPI2ZSHeZzT8MHqyJKPoYheODP3Zo3lV1+RfYZ/ZMeQg7
hG2xpQol1VCSZws+n6C1NjJ8lSUCiNcjPr9KD4b3Gpg7aVAj0Tf0KPOJne46wdEHmLcbhnbxZNDc
WNwVPd+f2ol26Gq1ExI8JOkky5NaHLPaBzC4zlDc4bVnSKKPWBebTh/jtcM1Y3IrrSTF5DXSBuqc
JCNlCIhQAjiGrPqXy30osY5RgwfSSkUeYlqnm70E7NJsn6G98o1KpQssAlrLsMkpG9nMLvujb1kX
tY1DQlVXBQfS6hkInwxF8kqB0D1ns8IixfbF3NKyTS1cIDWnxwksh1ZskwbG2HhInL8vFRBVCW7Z
kozzQvBTvNphmOIMhu5qTh0fXi6KFdgFZpRi+AapOoY099+DGgfacfd1DqcanVTj+xOIzrTBCSBc
NOF5KN2eIpCSrWnbGfsnBkLO0uczaczFabKsTE0pr9/dW9SdCatmdRAv3bgLM08qk+tf3PPq4q4O
RjlJHVOwjrhgBThiYMEaDffGsx0L6tb85WSMacbTQepKvC+PU9zlxVN0o3y+QbY4xHIr600FGrvJ
FqXA3pvIJ6LicQ2HLXOxMgDPFFjGcPvKwogQyCIpZyVWrN0FG0/Q8wxbBxhdxIC4fXxeyYVmk/0M
Z1gleEpAorHmDfr2NFns7sv1ah6PpedZXhLwXag0HAScu0mXOpNevaD4JPXIdGcBg7j8x4XlBmxw
NN777BHUXY2rg0s7qACcrkGjiI/pc7oCrX7R7baszw33dt2sx/o/ZIfuily21KQ+KbyLnwVi4c45
573VjC+xIWOdwGcD+WX/54xmi2AJgfzG37BX/MGmDYBSdDEc4sDfFJQMiPvwmNc4Fnpt4DPAaJ0E
paBitvVWJz3atlX4ckcwQayFoGGO7tp87f5D02mrruwZ5IlSKP3kHwpfxqX50sz10Rhl0ifmwupW
PNUAs6CNiGAg/zhE9z3iKQpEgWWVsG/psocVkbOyuctIcZW09ZVDV/fCXgSsE8VzPdA9f3sAEO7B
s8MGnv6oIGk5pvdNmgyJdvzTrJoHDy1yGPP1IPQ+8SRZHKPcs+BrwpGa/yhZPRqFQo+xM23WaetT
FxBqpiqaJpXzbILvSXECQaTWIgp0s+SQM2br4lEErSPHsMEa1aiWmCAlV9SnpsU2Y60Oiej22ObE
d70DD4nVyFvi2w0QoYAorFasdwuvo3icHNqbjN9oZw8R3Gowjqdb5jFgCqiBVfdNDoIFP0I0V03L
0e5Xp/Hful1sLiH0cNRi7/sFI7otNhA8lDX/zSlt5Dv2KfffhTwpm2uN3Xed2Xit/7YCvCMZ0lrf
ah3OV4X+UG+3oAdJ+bRs40FYzzYrcPQ97VkRsdit+R+OpcMlYPc/FhRwmClUp8hrm3elo4iBCHN3
y72qR8N7FkTtXDuoLLUghrJzxxX3QigsEKpKzDDIMFrri70eyQu8JmDY/2R9dt0jwbCPFHgGDQP4
TWIYI/vxwt5rtOXhFzHFkLGHMOJ5fs7BPeqRZix7JQQ2LGbqPjHjYwHHaxGQ6lE3GRfv5BwuTSEJ
ojLkYM2kbUjCNJL8muhEd25NdAPZ7TauQa3h4QgVYvJSe5uzOcklpzKzUbh/S1s3RnrEe7gW+cyN
zDHRAT6c6Dt5lL8/GWOZ1lFWX7qAhPMVzPZFHbn/UqwUV+0eBmxm1y0go/I0UtAqdEsUap/j3D+p
Zm1NFdF8KxhlUQx0/BEvbf5Hzh+ZHWDBKwp+FUyeONdpopqOouPaHPWdWRFM2pUC5bF3LTa5Lcjp
2RTVqRYJrjV/p6k57PsCuKbP5gSF3mxTpxhNG0ECuL7Sl4R4A5mpE3CZTMX3yRM5fHV9FebAsUi7
AQsL/iiJaTLzKz6LW1Nt9GTp2X3MQ1aBrTShqMyXVR7hjlUMamqmjSjdDNKFXRRFQhAQSXXVroxy
Rw9d/iu044CLvIEeG72VC6QbVjq85CaRL+8Me2VQ9hBygHibYMZRnrbqSHWMtlwmBwGNcNrxa/4u
0TCDPXrKFjZdo7oYN9ExF8+D0BCjSn1VVvjEkCTNCspShBcrbxJw5fUw7Px7D1Y8xkDdZGWv36Os
VYl2X5yrTQYFXdIEqe4/ZEthDuAE8WNYUH+ahOIpSXzuF3g4qgsU66ox8cbJp26PeiyzwHWCpODH
MZh5tVZWd5JE71o0n/9MMkMeR1Ue2XcDo/evKzIIBIfHxuTMjjiensxUoFx9AwQyiaTPgIeWLRws
hx++mdbsBqbER4KzC6xQJXb3gzhY0z5+3zE7ydXoYK5l0bCUK3fqsFkO+mwydLY5ZSmvFahmVjL/
warWPzaCkG4tv+XsbK/yZkytudJjjvHTBYL89eSLhz02RvqsYVJgI+ayCLmNxdk5+dGb/vrVsO24
G3xsdTSEseB82H6Opw0t6XCS0WJ3/sbHgNw5rl8XBQ5mQ/EPfyUxBgTTWBBNuOQTIDIFp3vQx1s0
jHLo+JUI3RbOYlKaFvOL7FBVT6b/iaPuUxDrkIzTLrqbl9yTvgY8LaDeNyOlieTZAv0SV5jOLPbM
zt0PSbiJGEc5N5ZEf0JmOPYT2MjMiJOa0GBXDTG6iz5UzAYHHHNJ8+RtrRWwwPNb/32YvpODPgpc
t1HZDkzcif7BFMOh4hLdqsk86Y5HRRZ84UuQZcKbeTe3kOrru6s6LCh0rdLyJ2IDwSSQF7ODrKm6
SXuggl10BilGn2gvDVzYek7lDlrYC3dmQISS4HMHe/OOLv2Wky+EPSsy11Z9RPXFdKA+wWZUF+z3
xoZUSRYZgFfG24JrQbak9FbGEcfs9j2isrUL6nW6zezInedJg5Vjb2p8Ms+R9GOSvNzUzVjXX+rg
vsokvjzpzA/GSW0+PiyJAC9/YLIESf6JbAH6qVOqxO1w4rnYjq6wwk81oqeIAxmxwMaNsXMHrusi
Q/UPCX4p4VnISTCF64yfSSV+1sOoRWVBrtTieKcEFrwbbjJyYgv+rMT0zsDJGH2JN6hO59QGXlEU
a7NZQqDQXb3XkONFUhQV9JVLUSrOj7mNtNg5dPRQGM0QUdmQa98bdiBIhtOK2ffeWQriVsJsLbdD
naXqJQOvErjnu8/plcdHqXn3PoNSUmFtOveMD9LjbfAh0FtWyVAbEGDPUT/fsZEcgHPZeii0yrT9
bdkKIBWJla+tRxr9jRbuUlhgfTFag0cE8kRtHav7SClsPGpWO3Pihn9nG9bPe99JPG7aXCl/QGP1
tDCCobChb0Sc5K2bHfsa+zjbCk//j1UwiLZe107aiiZ8gtnYh0BgSMOybkKgBEDnsDg9OC1DWbNX
RcbvIRJwg65yNpiKqKVWoD0jzvGZgFsvV707xKF9bbDaBcqd5hBfApN2wxx9q+7VZgSIlsK44BEg
+OHDDNecjVGu0GLUsHMi6JqgHaHJnHmrvDkbiGsO2XpJAxNySfwlPDjKpv7l21KZUSBNrtiAmBkN
zPmQHOixYwcVOOlVHxsH3obFCf5k87UHBwW8iqP6bcL8a+edYjkRtw0eHW1SrlQn3Ka45i6N3Gmk
PVLM++WCSBD0djBe+3M6eXCUo1jpjIYcbkVLMqIJz5iyNgsvwVbRNbqhkOf8AUTbuYfgfHLhjPv0
g8GoL5yZuP+xoLSh6OhaKk1ZFZCOXoJ+sCaOiGFqiKf8Nd5qHjCXHrSnuYp1l11mwYZLbB1/EzZA
e4h8ZUIryBK/2PNjQYwubaSbF9VaZAgd2KGXliokqB0m6ip1soZn9kHZKyfuSU8x9GpBW6dECY+m
DIIf4bgUMPwmaxzcuK5KqjdqA/JpCSGaBmrmGQdBG7onfW4gfqVn7qeMzOUv1mp6xryumP1NDGqL
DNvbMBn4jVQDxTP9HeuPNOVhqnHIQHamapsgLUHlvzAXcB8raXO8e3OI53/HRcPXyMj5dPt3Tadz
HiRSoCM2dqZsVhq8Ts0AyRXNy6vLMWP5kpYbquPESxOM4H03reCX07w2BCkP84v/RvGyZZMnrvua
Td7b/nHyj0v0K4dPXUm1k6l79NoJZsdC9+6DQZIELetbnML8xcuE6aOIjFzY6rtKegguuayFMI5o
ard+OlBUgXCYO8+3KsfVduRvKcFhgnwEisxu3Hc7crtZtKbqv54cUWE0SdtDBo1Ex8UPtdW+GgJL
DJmQjqLob1ib2qYzTXXvcnpdRi4GwzxLZ18hA1rsqUq9tcEGbBSaSe0poM7vOgkQvD2mbFXiGVkK
6kedhUcJCtARJ0bb0K1C6LCPkwdh4FvbkgNL5dL2mp4lzm/z32/l2BcdPL8aQ24Tz+Wvz1ptvSlF
hIIRsmdcon/kiugJJLQ4JqtW16AlqlesdtQdggHQlWnIXyH0On8hDATeazQ9RJrJvSBRuP1HEb5n
SVrIT13gsyar68Qj82RbrasxZ9Bh6yUZaBQfWATXIHYtpvVr2qiEnCngI8QavBSsPSlmCJsJWpJZ
VhXkxvtdNnGHxg6Tcmw7nyTD6jpgpb6sCgYhe5EJPdzIRfWkmRsaUn6PZ9wPfKCw/pZ9wpMJDA9J
ZiKpt6Zp2bUwpr67HWGuZizAqbF/2RBjRzYo5Qw4NhMIw+rHT2R3v7DZLusCbz1GlP/Mw/fr/dEA
MLpdUfH3lIHqJtiRkkjY6ej6X8nq5MT13LJwDyWTqJSW+FJr457Ceg/XZSbG+kI8RYudVGnyyMVa
HWVPUmonVKJJzMjigxQQkwjyVM8H/M80Yj0S8deEqK0lrfxZ6NjoaFDeaHW7z37ASClBIBNeVgws
xC2R6vmhFpN89fTWgMGdjLWIgQjNw7EdcBicd/37r2anZ3RfZoY4hb3SSeds1QJXfoWI8zxJgvWG
6WZM1NKffsXK7lIGVJrDelJ2b87vh4FTNytuf8BRibDRH4dNCUAIRcRYyWF4KUFx1nfVUFr3o8rE
RZHjbekApc8vMcTXI1B2elBfY0tYoxc97y8e1Z2M+QAjSn1uElpA4d4xs7/bcVmHTLKA2TLFBHTL
QN7fbJyO4B2zx4F4nGWjW2rlC6QMUHEDPp5ZV1zRXUhiu0+zx4e+pCidEtoztvHHMIhWxZIR40oF
d6QIg/b9CBqasbJXHbYIDCaoHX22H+JayEw4VElMc+z2Cda4Q3J0HwTlTDxQQKHLZrkbUarpjrDR
+Ezy98vWq6DzGassRMrE7rJybyKIyCH7yB7cSGew6/nQ9s6ldqqeTY8wUPyRc6UICKYAagPLdjKO
eJWUKMBbk62Qs3GsBAhL5Azlu0DyTJyVCiH/RcCXj8PoEhQOEJrhCn2wFVtMV8duoc7TKuT2gjIX
D/Fi7dieovx8vAtcFWum9aNx2I5EQe/74x7yIZWEZcx+XL3wr80pS4/sky0rMPR+kBEhPGdJXSaC
kKHAxdBMEncO27+9ls3+sGH/HP1Atw15TX6pJkHaUmtO2m83hNHAhgOV+8y/m0coZBduw0piu1Eg
Ma8qasXhk9kLdpQTKg3B249zEbPnGiy31oCWXiFnelgBFPR048A7qL2mzaQJ7bFd4pxJSVayXdhP
gYJt8OgmzPpfFE/k3eEhOVdlOKr4zz4tpyzpWULv2lJzV/xeHT8dyTccW6xeaMv6HU/trsN0qrhL
bpiCJLA/BaetWJuvyQqMheEnV3Zbf8kdjhf26/llA0a6uIXMVw7zhQ9FHu3eXjT96ETdoKCao9Fg
rra5s5c1l2fM6ctpWQsa1xPq4qtLfTXeD/emH3xVCuixtPyvfbN+IUXukdHft9Sb7svarPI+p3h/
4Bgmy7SgNKjMQsQilDA43sAEN8kKmzdBN0+jcGJH4JHFpnZFftNjOLg2P/5cmAv0pFyWpkTAnoaf
dJyIGWrhjQe5ZgZyfQRgNPe0JHWghlIqkr/s/BUY+mysrKdCsmTEPLd/drzf98S0+ukAA08/jrnN
qUXS2QQwEmV6YwNO3lQSq5YKQ3lWnIpRkxEF+eshK8VK1NaOFr/8rHO6neX7r1YtLK+Nkm81X9ou
yqNQjAXsFp45qOuPerolbmypW1PykeKAHaJcbWuQ3B6fKkwNESS23tUj+iUq4WDgbj5UcLoq5A3b
mPu6hbZat8/EHg+pVeUBVixCNGLg8yT9F2lQ0Eu4Cyfkbyo4pgvVjvrCD7eMWt7g33GdmU2anEnS
JG7FusHNrpQ/ALFy/L5dWYE6GOci2FikdlB3lWBfOIAxFSxRmzNX30Nah3PkwvzVrnzAnVvIRGNT
NXw8hF71EDRqWW1Cgtf0qp8C6sJSacn+T6E6FkAGb7svGG5IROEh6Sjh74Bi5a9G2GicAMCbUpuE
5dxyPFX6JsXXZ2GSV+QyDW3bvOdb1BuVmbxrhK0EqicR1AL3nOwcjmzGOpfiIkfvClgyX8TF8FMm
UD2PCtyVsfExXMqiQAqRS0Al2pracezjgS61J8MXGQOtr9OTBB5JGCuWvrEZkm68CGeszTrkcEbw
saqSQ4WDgqcpvbai2GJB4oaze9iMVuxs2WzwRWgv8md3mFum2Ch+hDDl1kCPHiy0bEYmfTOEXKWV
VYTOdc8VE6f0Twtk5Nz5rXg9/sPmJq4hjnlRDv6ASC47eCQXBlQ1/UWDswSSocOZTtylwdUESDTz
aBTqkXNHtGr9qN0tZEjF5OFST13JEvr46GQKZPSLTN13nIbZF0KzMj7GBuNMUubzeW5dMRVFIXva
b6F3ehYMX5bGzLaMcqKr70qbGA4g8xFmPppcBtymaHdlA7yjpuL/ZJ84FCyI/oWgtfn/QHDedECb
ITGRsPuTWWZMw1oeLTl/eUuedgHvp7FqyLlw6rsMKuByAD/bRU83LLojdYlMWpZ9ru1IzfIJ5Y6B
B80ofqQ++QkCnKkCnaTpDrBJtCXuhGM5TV+Os7BbmbzT0Uha1rF5OSBRoZwa6eQ17KR3K+AjYrY/
Xa77dZ2fsezBDYw/KzFYzBL290IHxivUmuwTXbuzMxWdB7t4MxrPSkGsMny/anknzCaOTELHwWCy
O7o1VDyJN3jzR1QK3PSImLQWkFJOWmqC3XxaruBhB2aiVRa5O2yHknX9dHmElYDboyUDllyDwRx1
i3j/YJkvv/xAYnTiMs0/jq6hJ/gN5edExxOznTMPyb68mOH7TJRjO/r5NWQLOvF0/JEgtKTO3zyV
bL/tmPIjDuwe4TrU7tGFwGycCJUN4FzVvQDfXVdMk5EaMVuc5GKf6bp1MaK4wUkcG/2LISOvvG3C
JS/IUUmIkyIkgGLDW1YsyKn7gmSvrp7tuTQLqv+rG4m5+kA+t9X8ROLHwy5IFF/9xcKHdnDGAGA1
bDMXA+QkbUqYXorZFpTXXHogl20NAdDDXmUcA0ncCF9acDRC8NwFSoYmGf4NuBmXJh1JXyWVG3mM
E7/cHsj0DyjO5nUoUyBvIl8D7xcOcraeE5h2AtA1pAAMHlSbA6ioFWM8zGmymwisHT/n+7OdF4kn
rsC5WHoO7Rz4KS77hcl11J9xqp2Gw1DCT+iA/78nZhLohxQ994J3RtqOft1S9ZhxkJjGIFxm+QPx
RQGfHiwHGvPX8pIuh2jH6mts1gU5j2XsULLiGpUIOOHxw6LR6anSIEczic5s87z5SVqFP35IJlER
VGRP4kKY6YFtVz/vcP7bWZX4TyVUq8n3nBaAfDTZR/vYG5pjGsoSHw1uB/ciRjH3JtVJF5432LWD
AVG9W9fxJVtQcl6RsREGSSeSztmRaB0P9V0v78gYL26wBVUHl+AzrscknJmy+pbd9kFttfbzsbww
sCc+NsQH385WYuwjOne4/Y9cYEXmg9cFreNz6RMzTtD/yM8JojDGMowX+t38WQsr0Kehzl+WjPqV
rvToUQy9HdTtVE8OsgEGeOOwC7/XzbbxnrRzOXbfzVyK+r6qUROH7d3/bUPzOQyRGXHVMj09wmwU
YEoYSzxppJMQFf3AgSvvMOk9xj5/d+j/Y4Yg6db/6HBYGMBxf8UK/N4lnmZ8H2iqDcE5cUGgkWTC
nJIZsenUEBYbViyKRJY5P4NwQvZmfBsB42rc9Hc+t09yMDIYYbiFWGE4iK7j1U+gyraxu5jMVi1m
qdVO5TSuYowLRZx164LQvgRhqnIEygcTXPf98/F86cRMmV0eDWozv+rnt1tw10JzWk9GaLdziRYI
Y/SLRmxspeFRKsPgxphcx7dHOZlfcoywkkj6GVknI85Vm2V4AwVaniNyymKxAw6jcXvBNuwpBjDy
Tyd5QGTenxtb9LK9SUcq6WharzJsagK7rqo7Ktu10vcOYTpgeNRB+QFl7uB5O+2fzJB3CyY9iExG
14j9t90BQFjAwOQiBltny1a1SBLSL/GSVDWzr1Pwo3MVO8LeAP9jkQcZzXSt8yGpBVO5heWFYQPV
ryP5Q3zjE4K8u7FobyPu1sBD01AZ/QWVKOsRqOif9fIiKynD5jxB7VhTPaLoUUKJouM7w27aC67N
+jukMBJhDBqkQ4xRgv7gZtqLmwXqW9s/JtJmUYR49kXUjX6L9cFijRJINU49WrqSgK47O0GCKDfG
/MF5XgBffATLuXbJeXc4S8TLnVr+RHOUUU6+sALfQf/bsJQCiBMSlR+zeBa+K7xgephTa/PZXKTN
QQDNiE4JIyvV+ffZqRRn9dDn/JvV7i824oiihkg6uCv42OBq5CtpfgkSxTeaI7W74B2Vx0VEw7Qh
LYDoeKmRvcKovgPoxoXQCzuMmw8H6gk0hzmIMAOp27SaVw+c6lOVNmu06Es7N7rjIfhuGBAvLRUj
iL2vzPbzfNcuectN/Sn72J4gtEiTZZMVQ3qzHVzbbMf5rKU56mvwVOna/mccQVPoFAXqDMsLbI0/
v8tT805ZLAM4Fr1Xu5rmeGcp5OtaEDn5uJUhBfvrJQ2AOw4g3FPLJGdBfnRR4VE6FZ3UhjSFNH6r
iMLoeMKaMqciFHR+UlrxSKhA+zWWvt+RTfiwDloZdc8B8Kgv1GVk52qyZWzMyfx5EOOMCzxg7C4Y
+AXGhj/+De5KA0r7322tcel3mwRPlxFK7A7RlqYd2B00PdzZIxE7OzjnDPX2omEd3U7/sH3c17hk
YkXYvR+U+e6g6WyGtK5BrHCenr05RmhURJWPs5fS4Q/J5CJLz1abNLDvGxVJMK/nG02KCzL19+Kf
weHWTyO8ROtSAzkSPegTFFqoLUiJENke9X9LuP15cEYXiaMOZwcMNDSbNnOm+uDCyXRmq6DBiJUw
mvKWhnikqh64/AbenBrOFRV5h8h+JdHDZFLcpK3+xX4NBFTDN04eQkC8zbQIOc4pklSetvgt6eKS
5n5p3h/8p0dVqkbWtbkfog9N1ATwZR53OM785W8x0vQ55PpFsotcIiP0BbXE50fZIkrDbftFd2Ur
ksDCpdxi0zWRgU+jToHGNbfJXqMHYP0zcOdFvLCuK+wklKJDadCA7rhUOUm7f3suzc4v4GofOzKQ
mRPAWcGLVuwSMmVdxZNkHYJMzXD40sSoDI4LaD5UFnW9e5XF3Lu/SZnTbaxhPnJioCRxsQ55/4PI
8pGvMhrE9GeTyj+Jag/0brusF7u/z4CmmQeU9VW2616KbijhaCFTueoHSoROA/8V/C+gQ7Nz10yI
e7BnxOEEKrQ80IHwGItlUTeE+i7b9MJAjBVDEyo9lBR2RFXy5yyONB2RPdtYZY+QxRv2jYOnlSrw
5PUdN+eHwt1hK6YEnZmJg3eug7TQG9Gu7wdGsdYInqL5l1Bvucb9dqRz6npV9LQNViahy4QFrLLN
GV6dMc5SOcLr2piCEbdnVYEi6lGVig0oRcyJdw8ZZfw3EoCpe664xOPoPaXBAJnnLF3NjKVUdAoc
3dj77vn2NvL2AGUkpSRPhjqWdgfIm7n73pWqOA2RVuzVddlHKxyKIDOpCxikc9KZSnhbxAMQ0/ou
8Ma2aBwmQAxZyuIugeAqezfHd+UwFOOasj/RyLSkJCwXgmnLARv7xXTKmackWrrpmXRY/pSZYRJc
UEt9/TXg49Xz0PZQOOif/t1Y66aQ29Y0zAQfg1wUVmx7Q1m3wc2Z8zaDgnDhILRpVckG6LOP8CG5
FGesL89s6Rf4sIjgkITiLSJ8bxkaOGvLMgxpTKXf6FWZP4OLIwQxM3yAKawzD+VlW2N/4jJvI4SH
bGYlUU/80oeEXtbSMMZEHAkrRyWxKFqM72XP1XDuH3x1+wWLsiYoOWkWLdAA1I3jzwa5qFvx4z0O
d25enSK/Ej03dVSrtl1EsQi6+pqa4Q3PHfhvbCUfC6P7H01oWtHkr9q18Kq92CilAAoKtNN+iWlu
JSMajb+wHnGMsg/rhCDKDcV1aFoOp/ePGDByjfhWiRaqtcvoscLXj+n+pG7JKcZ6ntx11vxxHpRB
nRan8g1Ow0B3solANpov3PIy4NlUiPDUAhpdi02lKQncDMc9FtePbNTxVDcKQkTXwjIqY6qOBKAh
LaJXVmyFPCrKxmwW708hIiC3ISRYvVMqV70vi6V0qF/h4ODue5wxlOkYX561LxwEkcFjQn/QqLlG
Qg3LHcaZjnOjdLT+gl1BjgV2o5n4ga62BuP4i40u+nakURSaRiJqnp12M4YEfrzxYkxevybWbsl9
gdb7e8zZ1veDKrF3Hl6ulgwJZ1dhiMeD71Uc3kW+J0kV6SlEuZJXfu+InzuP97WKMm9CDddUxweb
VV3VM09bHJyEaF9hDJH6+j2Cxc8dsIALDyorrORmwNo3dCPDFuFaBtswMNr7ZBAiIctiPVZg4O6i
S7YCORKxSDX1fkI65YbFY7czeTwn+0lz5KgJ9IT5nvDgo1xvODVpCbidlnEs4abnTfsywed/A7h7
NR9qOPcRnGCK1ZbX+2iu3mgzYozliZ+TUhFwwYBH1MnqLkdV/PsL3fpgvt1zCFTWeA==
`protect end_protected
