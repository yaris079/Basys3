`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CtRPLOKOQ1xvKzeLGjtL4WeMkpx4zAlhRzEHmyRYB5gRNYk6TihgjeCBs30gg65J5DWYFMnxVkW8
/vC2BgbNPw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
d/8fT4FgbYfKxMBbeWPR/ja1YxbO8YM+F7OxHD5BTokw677Ob3D7mlDOsHT8I8vWsgizD5bvSnms
BiPcwW/IOv/WNu3RC5EbJQthJlIRETJS4nQwh9KQe9DnsruG7YmF9NZ3Do8C9/0nc7ZcO5KeeBIZ
aaytjRkugvK3DCa1XEU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pUibZuP7z9gaelvMEZvg3JlNsuENxjoPiGpbyqPiRe5IHn9zRbY4EQdifKuGX2v+mFGYz1cTlhfq
bGuayOMrbmU6y6q+VNUeeYMnzWR8wrt/d9su4xhZwGoFa7GPbCgXHDYhmyPojkFU0ZUPCfn0mQ39
3o7XGY6DnyyGD3jzpS+W90UnuQaPoiXHRhbygZzSXpnCXmSie8Jva5CbtLiun91kNTclDY7k1DO2
IiQiytPOQb6W9wK5tdjHaLOquM+ap7l14+V6YWRu2+D1J+cZoKBqNNkGwed/hQb5VJOh58Pc5Wae
p6+IShXl6JzF93+q/1PUF0mKjBN7z2TxQhxOTw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
F/ipZ7ynN4i/yPWaPJtMNU3xCsT9qU9YKW6DApeLbE6HCjyVrCNWHNCM4atPwxVA2EwAg+V7G4OP
thlLv0nLHXbINEAO3WqgtsQC18o53EnPywrJpTYlg58Lig3TazGanOft3voJbEPBc++DJZXXjhFd
uCgG1gdbUK5IxpA+Fp0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
HyCAqBU6tZEM+VNYfOsM3UDsHAHa2LkRjXqPl7O9uTfo9LZKy4ly/VDZ1uCe7ipjlK9xL86ZPI/t
w5aBvBfJSJaqY+EVRjDbRcmgpwjIN+fSaP3C20MAiZmFTLcrHhAcyGjPmsQC4vosHxEJ+z+Q85QG
z9aFpV33Brl0Cj45c9JKThDw2s7yVpL3YUskA/WFISCGI8WJAKe+YuNkPl6a2JR+Zy3E4nN3C/5D
Usb/iuksxh89QwGbx6J7eEaGLr95B9r7OWi/j/quNw606TwkNH9Yas1Eb3KvGWoTkxicu3Njg9y4
xwvJeOq+G4d//cXzj14QLfwgW5mQyHRlQihNRQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5232)
`protect data_block
YhU2sESsVGWEd7iIa5mJrhc0FemyIxFMstutgM0bslpkksN1CHSSq7uh5uSJ3RChN9Pi98ws65o6
+cHh1sIloz0RUojBUdfGtmPejzkQzz1G2cuofz6hpYegWSE9BM8l8gD+oDp/07Ve4gqXci04LHV1
Yc4RBJoynNjKsSFOhot8OFEGvw5SWlhy4HQvDDnA3Rzja57kNc1c4jle1FEtY0/+jVdZXBudkKXy
4JQGuP3q88R3v7wwVQ+aleOXvewT6sqV8jtp6fY1StZd8upBJNDbBqT05SZk2UazkSpIGyXx7iV1
EeaxIN+/UAzzxHjdjrz7vSujNloMBCOAIX5obREIgvS8xcRuBuvWb3QpvPvDfB3g93fG2r4G6yJD
ATaCO5WPDoi9mzt3LqOw+fS9BSuEp3pB6FWTWpY+ggTQfkapagqeB5Acd1R/E/d8p+3QQUNSoKxp
1OGUDCbxtS/5JPaEle7OuQbZL9D223tBEN4T432PLI0pQ2gGeGnbwNMEChCX/Ibj/oxkW+YgTw/y
UULlvvP2GKo0JMSyXvWI5yIKQdRybmE4BtUpcHRJtLL06463fg/3DqoAFKvWWvNu0VdVco+cM7d+
3wKSjk1tReZLuu1dRM7f3wgAMch9Rmq6rYcU1c+RhJ6UsV6++UdIbOm6B9ZxPoSzM/k1VXVPZMfs
D4gfhsBH/4in0UHCSEefORaPPJUHCf5vhH1mRqH2fSdUld6pK4XYju2V1fvIL5s2HQFXnAL5+jH4
75yjuinzB1Pk9x/pzRuaAHRNeWAGEGDyIspo4v93I7psR7iN6PaMtgoH9/qeSz22rV2fVEpXFU6f
5XRJJ8LYU5Pkq9/67V2PZaNWMxKYXiRErrKg3fMT3dEmPJ7A0fhJolIt6haSD/6mxf6gSMVVNAmT
GcNvov7IRZCE6LuKegT81SB0eA649RFFzXyyWecCo1VLKcQpAEAckHQ0B/JdCSiACN/+YP16v4lo
L89yorv0DqVirDgZHPGyowtb5RiuyEdxjY/FKbZZBfSduTczxYb8ORa9GDpHG4IALr27tD74u2bj
5gOh+cZWarQJjZyqkT9hecoT1Y/B0XjDITCJxbFueOh5168Lw6JLFDxR/H+Q+l6onovdtnU5cwOY
DWz4M1MA7A+KsQGZ9ThAQjjovzw4yHk5fAm9cwacBkzxVggnrczoRthIdU5jtqyHdRE84emmQEIg
XWJKMS5ReoKUQf2Qvb6ThebZxGmC9RtPGKhQEv5++zE63toeT2leo2STHpp0I739c6aTSAArqLN0
1Q7KmS1YciuQme2R/1MxdYYKKvtd4x5Z79Hz8vWbruquz1Bw1ilJrLK6ht1pa3x5GeV0+DJXk1x9
Ao00H4X7xoPPLyUPPLatFsudExfYbZL6DvgVIk20Lac0ZTKWb75mf4uUKdCn1dwj9Q9DZelDHVkK
bt39R4ygOM0sHeVwrBAPnKrVPz/4SPFou8tMQlfouDJPneqa15cZHfJpqZ1aMyCX4iuNt/3FRjbR
t/9umzYpFLDneAxAZoUK5oRjGqFWgiKNEcK2uTcGwc5LYWIugKzq5Hk7PEgSPwh6osI1menXRihH
4m3v0bmopfbHSRLSVs5Ew9xCo3mw3dd+e6qFZCTpzHpNxusiI9/HVr82tvYNYrNYAga6zhySkBma
iGbMDSNA8AExm4wmX7mCM02QcW2kMG9dXZG/ucjYkUkv24N+FaUaOY5y7eJoWJhnisBJ3rAvEGf8
2SynnmKJpG4+f+TRZHY3MHzinFovR2I9QjwHWswFiCKusyuwCXQ0snsFSlT3GyuVxFkOJ6oFJ9c1
asmNNkE4zH86Z1eBGV3gbyXUl52q/YUt+u46wGGkSAjB/lnDJlCJCwIo5XDFTmAae0FpTGiaf0py
GgrpbzHu/nyC4W2hkjr6bCUV/YtZA0G7viU7KtdHfm4j4q2udZPZ69MTpYiCeciTlk/VO/GM0eGp
sQa65nC74e9bY3Yj9Z2dxrRC4/0cLvnQYHDXU5JrbGz3QxhJazFb10UYnHExgUfS0C+veyOUySuR
xGnXu28wRhO5iQyxahyi6HNGUPBgX7iK39ugdA5tI/h8Ub0KrQe5UwIVAzmCAt1c8QmlZhc2F9RM
H7Es5+PUiJOL8P4NWnoM1xJtEDfkOcbIGwVVyVT28VcCoNFYqBNj3p6z7eZL63j5W3tKe/6a/tXG
1DIAOHHYmcVY9OVlONIFKz3XDSy2Cy2yUebYd09PxfJZ0TgkpxyKODI7k+1l7+pT3s4YX+6cCE5o
DAGgdzdAPqBpAHG0SxVLGNxHrmPKQFqXdkhkYOkjQloj/OLQA3U8perksM8lhO2Gog7zoZrCG0AK
k44m5qCUVKw5I8uk5tddeBbCN+k/Q+OfJ416pLFq97w+ViON9i7/d0o96ZlnDmzWQ1RkpGQ5Q02D
d98kDD/NSz/PZagqFO5K27L+EV7q/ZjbV+oMvg9cLdY3Gg4twp6jdDeifdO+FTOtM0dWqN7WSOWz
PdR7BlliGWA4xO5NqiPgUFLBhQpf3hVOpZqWlVRkClqzA11pLh/OvGIsSFgozQWh5xqRvbhFFTEp
NdHfDA4wkQp1f7eG1ZhtBM89QHK36DQLuEbFJZBo18vXkx5HL+y43bStF1zCSX5sGgAERexNxjDS
Ua8GUpjNHLc81N7Lmu4NEpKl2h/ZUHkRJHZrUOkU8jmerMdstAWIYuxcgmNCqfLVleheL0j7IXBF
J4f9zos05MjtjP1/XOrCnVMxMEjggg+IraPuuvJepmxB+ls9X+bLV/5b6r+kNvJBR3+PTc6KPlTH
ocQ95vqEBf5NQ/Em9/4RX3zP2RoMy8HTA8SgEP3XZasAc7y7FUpwkgywEBlWhbnMJhs+lQQhS2Um
5TSp9jP7aINoSCFxbzRCEWzboxcW7x0zlP0vHGixOoXQBj8C9CH3UsexTL1JBrXp9jbxzH3v9RMP
u74GJ7FWwb1CEgHwZc2fIl3AFf1Z9+EHXzW+QZbClsy/U2w7gfXlQ2hD6+83DbuzqszUtQiyedw0
fhxsn8uA0LcpO5yakhZOA/snHcvT+Wjo01B5xe2xEEhnhRl7HFO1oRtooLPuAUhVyWQNN0tZG0e4
VnRHqHpPWIRz5LcNlO1NTNaSa8iJ8aI2027CZaMFaQSfIXD/tWl4/C23nok1CF9LDDAGete0SeMb
eynGcaIIb0KS5jeo8q7ufe1rjeE4s9JYL92cI8ED2bvhzsobJkAFSO490KQ9x6bJ2rUle/n4op3M
dqiREpRnfNAcYImk465LRlJ67oo8lMDKC5uLSi99XiGcndncC6I8+mss7qZ2xoQp4s3yjY1fT6nJ
eW0F3THjn9VshDLgVjek62kFqh/wJ7uK3qc6AK4ZvXhn5lED+27dpK3hNXmYWAQC74OUU+fIhkd2
5MN67P5arw9DPcfoP6yYoPpWp03bImrvFgUsQd/FP2XOC3UIa+B3FRR/EfbZ2rwKlaVNr4cepzm6
aXx6CRymIOYt0UxIXeuV1MBIf0YvljBUx+Q8REabyAKVxLEeHIWVy9wpCK4EGNKo1O0Z+VTnz7cB
lQ4srRBln3hBPbnWK2sZwxzJ6vX9T/j2WpzStd0xMT0ZVVb0T3EwrpEIIYZYJJ+lvavN9zmlNZ4U
HbgrswdL52i5GN/DkBcoJc/KNI3RhVYcydUV4FjSfBPVdft0l68tZ15zR+QWCGwMbc5MS01xS3HO
oyeV21fDTQRdADD8CNAxGW/F0OC+CJg1C/77haj0eALk+b/G/4F4fmAPn6k0ei6YqAROeat0XfX9
BICcIwMsRcwDP1YFOhJ9caGA6Q8cYb2pbl2RHTrZIY/2KgtDO2GWq58KGNYfMXkcPJn6wQbr6RCS
GKRR9UG1gbMF+oj68ACxUO08b79ul4FOp/fDQRFN+SIB+EDOW/5k2Pb40GI1hvr82tVrCKe9k7T2
+GEQSad8zmaIgipaAOZU4pR3lNy2mBWLsbSK+8Y+VUs5zNIaYw7ttA/TRxp4oIaDFfR/Ztxeo3Zn
oC6VqruZCX8Evnza/4TXxHhwITLUOpxCDY8NfgghGk2o/7Gu0/RAPunJf4Qxxo2QDyrv3r1tvicb
n0s4BLZPQXUTBw0vZAZy3OEzKLNvHBvtIInjtioQgC6NDvj6/Q9v3jBkeV9brXst1CsAxPfN9tPQ
TxRqVd5/MtEMPOwQBLOx/I5iL7amzVWmDLV1I5UvsBmQ8rReoclTJDWFuqdjXfZdSu4/pLC0WsiW
tCTPusx9w8Oox7M0xx5fHNpWwVcd1FYEC+GPT7S92Eyux/HziQ7L4ZDWlVEcg0ObvNELXrlWhawj
dFVQc4MPyQuYvqr9Qlljw4kFijBuIm+Qwono8rcU8hZw4RMg4rhIb4pQKmwb0tqamPRACOhmbP2r
iC0OQAPKOEc+AYymFFAmmsWAgHAYx1qhhp1GMdzFo8eaRqOuRgNPmjfMCaCbQm0I2FG3BmdtsXxR
NxClgsubdUEirWYKYydzH1zvBUf1R4MmqmoOmFIC8CwHaj2RP0xNKi7EvMrkGf2VBdheuchIH/pw
3+lqgrFUcBFlA0TO+OdSAfK19rSEE0jzPTBqS8YhzkqZBOc+1IMU2OGkEtkbHNIjXvRZ9sInQehs
4gcXIYC9zV+exDzYdlbmNHZzRxQgFOaaaJS1RdBq7AVvHMHYdFUot7JjDpztkWDCs4cE/uUU2qVq
k0JsSv62iQohXjnrIknMU1TbUopQg4LBOrqbdBUYGbop0lUfUirST1dy7PQ/CzcC+6ik7Un/LKdc
8hxxnku/3Fb44kf4VnVvAmu1yspPoq7o6GRcRVVmkIZEySRmu6JpNrlZ2Y6AvnwGiOWA4xQL0XRK
R0NosZQqPYlGRjzfI53NhhlfDZAaxmy2CvyrzgQeclJyE2/8wFPX9yEHSajqcarWafAKUQbFGYO/
EJX4UHrHcsCYQ+kSXwkTHiW6sb1EE0h4lHOKeoTlaxeGS5qE4DZhSjEFZrVRFl1HHrCjkD5AHWM4
mNJphj/XjlLQBcq6frP8PR9DUpfvU5R9x7HZy1VpT2vLKCcZl7Nc39EPZ5HcX3YAY2pyEXEDBAvs
L4/hDgBYEXGUw9By2NS8YJWsznsB2WlEtsHm2QpglJdWwbD1qU5oSaaqUmUI1jgNE8DL6ihqh4cp
kOhEIZRrUVR6gI5c3XiiEC+YEZDEnyNdHxZQepEL0+51BwcmeL1trWr0AKCJvzY8mK6KeRHCA0T5
eAA5Jb0Y+crk+VfZZIxAxINypz3qqSfb0kKpVY5EyVeOoV2cCegMsqHFr2YUgYwWH+N9robcg1cN
Hzh+NVp4V8QsDalJ8TChBJziYlgkkPahXu9KgpxiNbK7Xt3LUe2wU23X4bTySoNhBtrjFYP/nJEa
H9y9rKtNhcsGsVnCvCejJ46/ugb3vASq5GyzqIpwnJAyOv3svA3ElOhIqtqhTiC0BjIVj3YH7nw3
cFOLzC5zt934QdRfopzwuW5wpaxYDxQ1NN4iBrys9mWS/TGpPiAd5IyST9kwi9Qpga13vK+uQg75
oA+/Vps+a+dRm4gxhGbP1pecWJFl+N8y+hREOtZzslXeh9u/07V1h/KXSxR+IPRHGSGQX3PlF6jW
u+bWN1//UMQOjAhNb1oxPwCJKt2fZSUAPhpaPfy3KjrqMy2LB2JIfVSs3bOBj0dk339YcikbeLzp
UUG2Yd71LA5j/TnpGRKu/M1av2lwfw8GyAUJPhqY/ntpa80SHsk3iUhorBPbhYGql7nxMmfvUPxK
gLYPBI7mLLACvXBci8fvZtaheaDUY7e4bEpLEf2RkV6Ije5TA8drD0spHkhPG6kDBwJqTTwYfP+2
a0yzcekYmH1e+gAdFY0Q5qV1PEaoD9entIQ9XCQlEmZVn84Er24E4xK65WXUgPlnnglqsKLaxYdb
ugxo5JIB7ckxCg8UZH1vrUDKutCOGwSXuokOb6f142oL5Ozgiq6iok2S3CVr5H9yeC8be45YhLmi
UnmhWLYq2HPjWitxm2zmPqqyjjDm5eYZvKc387cM2odfiadSPXpvhAk7QsqJXTXwMKPNRYDyso5o
cadwAF94epW8mdC+7DOKCWeV0vk0i3D1oJBLOhvF3CKM7q0gN7/v4R5NEyBIG3NdgmyYIQqHhmiF
pQo/0FCEbOKAMGbhVAmE4lnwsutJXFpDBBhovLOr5iLsCMruKClianHpKU/4l4N+4P8YepJDOteX
f8VQaFoL8mX7UBBJ2gJuLjIomundgxst2M+UP81WQSzW7a94xmDBFFCe3frazKs4Kv/YOYWVYwy0
t5PoYQZ23zoBFRDYCQPQiPJxSol1FFCsW9URUAjwZ///zx52NzH731bXlNpvnZS2P7UICh0vpm2j
XBd711E6Z4uVMT0zdhuCT8ybBjSAFqfcZMgcasMPudnHGVjn+WAG8QpD+OI/D8tnzA2tMYzMx70B
b9ibNHqX7IZWzklQ6jVbpXTLxVZ3Ip67cmEYI0qj4CV9XBufhfywlmD+vAv3H8V26pVML9wW2RPa
J2+1O669OuBcmKX5QpjzdKutaVD/HXIHrazueLPq4cAdk96+fvSuskyYtuaI9BisEZtHlVuUAMOV
s+/gO/3wYMWuciH6JZIHI2m9COQUMIg4ha0vOMW1jx1Ks3/ZogW0ocjPu9IfY8ltAwxSsyIaLgrm
5bw5LdCMF0RDRVJUGw7poDqhEEjqU/unte84u0dKAFdoW+9nvhpcAnoMp6W4HMl/wbqeqAfVDu+N
YoK1SK3NlP5FOMrhdVSWnciqAeEgQrC1OARPY2vZHY+74n8H4gzfnpDEl8DLvYq1QpFyxV5dMwjA
zJ822zZJofCpHagthGwsV3QeFaJdnOLj3wSTnbLZh6mutC8tQdBrgvc+9J86lZZ5wRosXDfYtuOM
rLZi9D1R9kFRMPdtFdvldV7f7MMU8dG3QZsJ4s8BOQJAJ+X5yeLL4WkybBHP
`protect end_protected
