`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
bre8m3ch/VFYLf4pqUTJ8db0MnF6ddmc3mKHu8iXsD2PJj6dLZdHWhJ1zBsd8rJH9DLMN5ebPi7E
Nu4TD+FtvQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
odIem+nTBDzlPckIHS5HBsSq8ca0XWfxhv02rmJBL7kfh/HDuCKSXJYbbBKxIcGiEtPlu6IFnsWu
2/CVS+uw2z9JTIx/w0A5D4S3eIVHKD0y0dSbHTXYVLigOc1ZW2bd9qGXuvg6sr8dBh00LD1hDuth
rfKIvM1tGVOBPT7zAcQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
W7E/w3iZyBtgU8z7+Anh9C2/NfMOXSvLPLEVI9TfwINsFYedcgETla0kbg9IFvCLoGYyld2Bn9zn
et6UqJnseuLqCPsVZq/dqq7CiIDTPVaD4X5P9pRB8W/ympaHggDUfZjk2O0aHwnDRpc//XuKNF5Y
wCU9UPsI+lyZ9SRpZ2iT/CK1KLU8dzgWotPb6BCztZg4hTXFAglfL30PszWpTe9ws8ITv9jgLJna
Yk3ICToRkvVN+UK773ugOliy1IX36cXoizou+eUQhSkCpUVyLAXzYQbHTsVfo812UIBU04/keXd8
H94w/Q/Fh5UK6SQf8IO8rovo83eNJQvqnWEMAA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fEpQD1sSl/hK5QTT8zcWHuyLVbpa729p9DyW+3dJ6lxS5zTDiIT9gWIYJPGkOj/RBJQpwo7Ncr1n
E/WnIKFviJREe2RG8Z5+Mi33kqV8klV0i+KgXy/wZ9I7ww1gYLKNmtRwQklzYDCZ8d6E/uD+yemA
TE0EqFcPw2020j4hvK8=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ELBuJnJ2gk6/zsYn2x3rzW5A40KhjjQBQbaHb+easD8yd8Plcs8A6pb5k7XJ5/jcVag7xBr60dyg
trVEskWlf39A3Sdj4Z5T9nm1k6JDvHwY/NF6hk8zqGB8Lf3jpxXhzTi+de7t9OqTtIlZoZXXXrqs
nOVbT4jgD80/SSMeuH9wl+gauJoK17SSX8D602zuiIxTFSsnxx5CzJPUIdJC9aDchXF7rzBrdsvF
SdrtRNlV5eBiZy8d9YCOiRIa5blzd6dcjPp82D3qYn5qySZNEhZqgz0XBT4sHsWmS7NsESdWutQP
WgewAVT5Zsx4roYCT0/EwMFFbl+loPvj846gAw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 98272)
`protect data_block
Agz6RvIsLwoJ+2SfzCKD3CiXL19VXSpmKjirfMaU5VSjdX+6WfnDZ4Zwf1DbArdlyBozTfeKtYkf
GB0Vl/+vr1awnjpZb9R9YiuPvLlM4Sn7sN0PBQNHecMzvhbf6+kHZuhJClLU1CR3jb7E64mGm/T3
OD07DPufocv/wP/HLfewIGQdHIVn/by0VNFVKfaqkNrpPpg9nabunFXydw5s6DlDjxg/iXQwXT/u
VeOdS2M9mVGE7D8m/J7ZNrMmEX1y3I1247gX1rQ1RxghfobQi+nLj1uAbuvOhPjRfu9acRqXqRoz
ehTlnGacVpSlqtb2Mu9r2LeZ46eadgazXOxW58VfNKAJ0AX7ibBjMprD2qIlefzw4MEMeeZldh0Y
1hbRRBS303nE2eLKfW/ntY5T+3z/Bgd3CAB+9M4sEtmFkUe/cUv40EiC71WJs6Mi254vFsmYg6vI
Zsz7ZvXQXqP4UnNSBlDeooJy7uRr7Ky7v9lrIJSSDrywzq+83PCSnv5pH6LSR2+AX/XuHcvq3DnS
vKhgj0vz/tSAYYLvnVBELQqePrAfFN2spiMUA8ipnTaUuiURnKec2dBQGWtgqXsD07dKy/Klk5rN
PCrDJJZk29ymXUueoEjjWPyxKG/spRfVzCUZmAvsPsNOB7gzks/+TwezgI91zrVCmi+BIYKQkTXN
NKH1+c1sH2S7wpNih4bONiSnE1d7+GJ0BmnAbWRokKeBzvsLjE0ZsBgMqrGgon/tIpXexXPDQL7D
G0d1I7okmVQuoPh4vGTqL7tzHYP4pTPn5JzgJ3ViTueg+FTmKufGi9d8SWNGbhn3sL4kNjGJ92sB
fmBC4EfWlGqEYGet0yEpp+owoWK92mb5dgDKTlJsIwtnLGMdgTbEsvW11Fr3OEoq1toSzgalz2hv
7/fJmGCWQOjD56CmFHsBbQj6qSA0DRrIbeV7TULc6vZF/e4rLe8iEWmQtW0PJg1kPBrYr8ldMogL
Y/JHVIQFAK/k/UbxsWwafdGZyb4XhDKpeus4baHgE/k7ZHltnz5lX3EnN1Y7k2/cXyq7/XIovmP7
Al8Gyzhv7eD9h3XiDmT+emAal4bo9q/MhELzeKvgCLdlKGej+bVAALJbAWMDiNnkdTPg/ef7+AdZ
5TfRL4NzOLEJghrWNE4Wm9rcj9bojgzjlU/PEayO/CesjCYbv2LYnxvLxL5H3Adu9FGuIpk2uKWa
Wub59PGwwZmkTLcedqjXbnSZ7ZFC3AjFSWq9p5NFFa0X+3auiX+wjjh6cgsm1ogscRH4uH8GfVcw
uCEpCW3iJSHi8g13hDGWsb5BEgejEDv9nzXFT/KeW7ZXalUy83N/dseaJzMB+CXTO6Dk26IyzrJm
6IrZi4BsKOW+NpG/IAFEtiHwKKrOi469rb1IGz/oxMN4j+uMiJnq3DiNl596UYF8IJNgQ1YYeGvu
VLfmVtYDy26FBtnyHHqcQ/Ox0vs9jSCR8ahM51jI9YDhDD/3LuQ17SIhP2TycPeJfeAqjVJJDixM
zlTdO0oq1bjChG6cjgUU/H6MaWT3aSnuEOAp/Cj5as+VgSsPTckblCBlUmtNhqHcjiXPHO8JHdhH
K5CrJ0Wzldf6BuIptfWK1NEM7Y0uWzUj52ewSRszXxyZ2fuPNv1kDWAhOweAwajvMU58GsGYFMm0
1JgXo6EzMItq9XxrUl7Ij6GtCQ52jsDmYEra3r52Y254d1BWp/m75OWa9DprrKwQmt/H5M2nJcbU
8RUr9bEkIu3HYWQVvP6vakCt71LyLxLmK7GYj+jVvOwEgWOkJwlp9Hah/l14UVJO3LWDY/vGy0mU
i9hQ3lBHXOx5QzwcHEt11huCymoG5jEMAj/EyQaGai9LMAMTvDJZOFZuzjhBNWuB2fmC1dBZBvCg
BNsDmLSpWrX20F8Z85Zk1zvXLIZdCOpwvlc2KJl2y5sstoE6dX+GITjN7u/VvUvGti9xuMg/8DsY
5rtdHpq0YR9rhxFoqxocupo4cP2aU0odjpyXtua+RxxvFb4coav0GoatEdxM+Q1UjvVt++E2f0Na
QQPXi49eE+9ks6CpcCvBxuo2hWfLDT9dq8xYxLhXFWjwsxj3hMYnj9aw5FowljuQcE08/WmfsTeQ
5elm9kb6AmkRhHwEyyWJI7YTS9wdmO75of5Z17f+0KUQNDLez/CFPGL2YLd9sP29fKbXt+rIUIct
AnVNfwuaj1YFJdH/WAr+EHziYYHWtvyF4KFHg7xiV1Bbx990bgJf8pZGiJ8lMpXYwH6O7NYKWrnP
uJfLMnqCxsKrD8TIR/P4y+2zg4zlPvfQUh7KvqN4eA1GCFgXdcl/LjZfD4elEDxq/mABU3l/9zxm
1WbOsVybBUXYtXVHJdmud3IlrtZonUPRgyktWkJHcpDx17VEvp8NKtdd1mL3L4HVo2SUUgDSL+pb
yQM0PDJRaU+nox0MxQmhpeCXvCswtv1Bqa6pY0qGzvKlTkeIn+kzFHomP8cQZBPUifrD+jmpPjvE
HQTDIP/qBnOgMB6oEkIgeuTsZVUwYYJtKADrpx5mpZCW/ba9QvLp7RoaYwybjrMHNRajvEnlaWPG
rWl4WT4u2fqRtiGw0fKAnGCfpO2Lgxx4iKuI6cKBA5Y7TP4mQlP6X5V8RJkigQyn7rRfmrtYtEnE
/1zsuApT/SIbyQWLMFdJ3gLZ/byAkyBIToZi2KiTB/1a2onrxA/lEJYI786yPOEXR0IqORbMIxr/
STHLZjyYjuRBbNEeWQ2B9oylhdl9nlphMG9BY4yQMU7eU3eZtFsDvN6ZgpEVR77f6xYVZ4deVWlv
8QdMnBK2NFcT3AOnMS0MqGkkoYufV/5cy50aE17yb0oXeCs7h2ff+oRw4hAgq2Rj0MCA0/UxMRl0
Q7m/25S6NofqMBPy4Qjz+cXSw6Wl9ajheQxZMbfLZLGMAkrqE9oezD9P3HulKt73OihnXguuabL1
4yZE/FQvMDguVtsx9CaU78HgutXa3OAZgRM8a/D3QvSxGGeyaMvNTTguFMWu7TIbmKYMbcLEpchk
I54JaxAhQaELLJ1vznzYSVa4WIWtsukVq2SdqGfYq2I3FsB9ydRodSeUJYnsIzpWazGI/z4SLu7j
UDLc6Jpl08llh0+izuq5n79f6NiJ6KAyzfjl83cEiaGsHUUgUtpLwoV97SR0GMFr0Y0w4nx5qxdm
80NIjsakTERgjvcxX72c614bRTAJzcFyq06exYTgguCzo0Hi7kpjWzsZyQ9bX1GFUcjOp4epA5lx
DgU+d77XkujWzDPp02NllF+xSwqbPUh1OFxO0ihgZyJTk8rpSJpJnEUUAeKEoyfh7zfNyIjnz5db
pMeAnejufGQ6FbX68yJPq3SX4RoKBSC4rJJPROkAUvwgY7ld3991GWtsDcPU2Hz7I1ZU5ibe1XSl
gpMrlawT+4WvVW6pD+nDFbMcaVzh+LJ3EXf3c3239oMUlKv+S9WktKtMDQsTnHMvMwwq6/kzSlKE
YzXvPB/ONhz9jNO4mHBB1cLLhvyAD54qqbGiUnzWIl54n2SuF6MnPgXkUU4tQxPR9zrlHZqKcXZa
ZsCA/fojw0QT+sx4dDDFNMm8A9AsiOhzCoZ8VY8nahQOJm0v1YN7+qWmx+iNJypfVDQSV1Yc+A/X
QEil5+TVAHsuiGYqKTsfP4ekjfqTXzPxburIsu8uCiVDZ5emfroXyyCTnQ0gz7Rnb0u+nis1e+l8
4rneWOjAdojkIIVbfODef6ANp+T9NGy14HdlUwM0oxnx2uN8CV+wdHyMABcmpagdl+Y04PQ5a3jl
jxjAuiVx5DR0BeN2LehFla2nu4hLMJK0vS6BpAgZzSi4lkOsq4V84wA2j3CPhfjR7cbD7AuBmaRm
8Y1TeBAZnwj7VcPlZvmr6z4TzrKsxfXqtx8Dw4dlLjzakuzSo4mNF5+QXjfn7IGMu2nb/YsY/pnK
ghKsbw/ebrqM60kGP4i16jIrV8Y3mJJoTUNKoHzw3Ue9aYfoKJ0fNPFgzsANaTIDQjR6V0ykqKZZ
k+WWuj11VlenrW9zQLPG+nvpaScmbHHAWV6kussSAOswW0a/81Wdp25d9SoyiFPAclGsEw+xmINI
OCXkKJJ6BvzXGoZPRa5XxDF1FLaX/khdS28/GZz5LMsRyF9kDutD3z0oKpVwnGenIcL4uB/XzeR8
OjwK0MCyQzmGW1rcbS/TDpHJNRHC1+KclIRBpCdMRuX9gDJ1jI3LbrdXeSUlYDe1a2I7+WbYKWaf
vA7HX1nKLfCbKMDM5xK1AWjqa936iuZ///n0U4gAYWCC5YwghVHw3n+6RSmEx9dRrq/zQDOwa1tW
1IDiRDp+FpTjj/42H1a5rzmht52Nh4DPCdrOWnyteYHenz03VylhwZagBwmdqoQXB6K73nRO8vhF
oFgx1X5FX2WZluYz7QuDz46qgmXvq/iixaajYCHMjTh9EdBxzqcFQD1jfzUdZNx85RxNWicF5ABk
mwwxc9aelJJCUPpTm9slXduZ8vDT2TC6YB3Jn3e2kSyo4f6ybI58GULVI1y/LiH4r5fgcVf7AGe+
EsIrsRPrsRjHmOOEjrfv45A61RIdOEeJRtIsqCKj8YdFi962R3NppMhCaJGGHBRruAue1pJemYgq
LYehWc+E2kAfHEQzvNJqTMFl99M1r3MTQTlOdwvfm7DXLq8jDdRopJtcw4re/A8BVdezgV0dE6YC
g8/iT2BCkLyBTje92bnDPcIwOmJrNSkbTpQ2DWJGANE7TwReJRF3adExJcVQtO1VXVSJQLQmnnhj
JioHOKJNx07mzYfWaU4N/2pOUR2Ee7LIMxog8LvXeOdwBpqkoRVBS+jiS2FDI/umKG/csaFJll5g
mZp4vwK0m3k3XVqCeksAWPHhjm3LKNqIq5oEhJIT7qKqzzHyr44TeizcMu3AgIbCi8fptxxvA768
Z6ZxtkztNTtVXdOsm8x/Ww/mhjIv9lNQ+LHsEcxnnuy72AU8DfkfHVZ9tbjG7lhlK+KI0M9H25l1
1goNdfTRVzMVgd4mRxjL9Jm9m1l9sC1Fak3pl/BtNg0qfgTWMWMv3DMe31VjIcAk4uwb2MEvNmOx
gSSA7vUOnZVjCNwmf6/64f1e0iLZX5j+3asKgjKYj0mK19MydTC3BTZoZs6nGgPBHQzvBS/2rXuX
GgGw7OwBU+M7O/JDPpfyCEHH2fGi7NeEIxuuNlstmSKF7dL0CGbAXYxPDajb4WkoicDwFPL/3xhN
KMRXTPRMYLPLDP3g6BIRBuDb2EwZPGBHIac5r8KKpPxd1DraO+7kHRp9r2lXu02YZ+C7Dqn4ostx
6q11xTGvNVPJtgpim7BfRjcOEU6oDnm4bnguOzDPKE5J/19PGRPNTv98aLg/QaSV492ZNHos7oLa
bSJDQR3E03Q3jCWj00iymVUTlPGNSjbthSmRWdIuaWVCIlHHo6+Vj0/o9WwHRESr6BtyuL1ZoNBq
vhgWyNWPEXnGezIrpRmvm6hk8PIMff7GFTu3IyfKAPOfXpvsLLtXc3b7kJvU68ibIH9ZF2Qt65eb
lGUUIQ5jGKnarSp6z46RxNKQJVxDoBpPa2mea+KADZ4DJpPk26C8949yhKS5F9vge2jxoaW/C9P6
NDJCQ4Dr+gZn4gELoSNkG/BJ5g3kmCo9O9ZGDnlt13kPCt+rx/mIrM/oSSGq5ZpxmOyMA7Ae+WFg
/7OV9oq6nRxye8FTY8F9ciirBUTeg5RFUlk3Ao6h8IpuZRslCxnq/ZwHd/cGda+b1jBo1SyEUVDn
1sRfVvWC0VXNhAa1yTYDnXO2yhoXsjGEAv7hvEe/WDxboGy07oAuybukeHYS7ebQQbtrPEUP21ko
KqVzKuG2tBZQqQQW542PsEifedL4mn0OpiDzF0s7LYZoGdcibV9DjilQxP0j3MWii5cS6LUm9iIq
w5HFn/aa/56uCFF9ixGN1qVVjQWMYvrRZ+qJIqOQFMgBvDwObsqWopU0OJlocAOhddN9vpZrWh5l
E2fgsSrhVsaj0q+DWbDl85CwkEC5B9KgwhswSsqfuDd7kcupSaCNPJh4zN8w9kPm1ZjGbNgwW8Xh
PplGwD1sAg1UST5m6SGKn8/ZibKlsf+0rHrX+eQ+EY+xixwR6K3N6NjBEvwqRzybws5TUVU9o4Jq
KdyEmAiftLAQCYRs21EEahmDb6K9YK8RojpqjhjfT0BA8lp4vbzShZeaWurjVgIT+5zgqqBsMZn6
4Rpo9Z34fTfdfJwYZ01RZSvK9le5ZVQxqDTI67L71xaSeHjlJcteCZwNGa+DOU8xoFxFtD73nJZp
SZn1GKUD+tEREzVF+rKp2lCasjmXEVYrhl14jBUZKENIBMYvnfCgzRrq+AxuDH6ljZxbPU4qqCPY
xCyOXLBhVopBGxbQmS8sfmzK9/x6uOqEXZ12lexDKPwYL4r2PTJXmpWx7wu704rBvqR8/IuPK5lP
TsgPQc2oy7BI8d0bKy9WqAsTqR/iioZ4l++2yA80rr9bFRe5AbS/3y/qwol8m4Sk7IHYweZhpVvE
VGVIPCBYA3Wo7aRBbZf4Fb49jw6HTqvnZfSALFVeTIAtJwy6Zw7uINqkXRnxXLg3PRADlshQQKdZ
ybpLoI7FFadSsl79n5fanwalRR8h6vehoepvewUtkmUEk96F04PmHxXU5DKqox1c7SLglwrxI4oq
dn25gWZ6lxZv/vZxccNhe4bETnFJxxbabQZo7nyqv13XnZY9jm+3wCgkgWGBJAS/wnn+BiDwGYKR
liPtaE/x6deCjV4YCzAb8OL44RNwWUI03d1L3OAW+IQnA/s/YbAvdxWQnFnxzFuUK/IBDX/2Z0QJ
lqp+yHRm5lpD6M8JibIem9jneNLhZCXo+BVusdwb6W15W3v8qwzV8CXOMMgzioJy5C5g+zSYZ7Cx
U0X65AA0evkIZ6TE+G7c3xz3zCihyxwr8amb+r/ztfBOYChFl3OzJXfxz1l/qlZF5XJz/fyj6+T+
Zv/v7S4Okq9JhpJEphUEqX5lwpbrWwzOJHpTyk25n+3tdPzc9097DRAeFZv+pgQI3vDAXp84EAWu
qxzVe002qUKPLZ0FUgesHgosjUgXAQG4jUY/UKahTd42gXPBUNK4uA0kNjtWLVeiqbOVhvDtDA7F
QMi0CEftAMFF5edar0pboFewwsIM3KXvB5H3swSIeJchrZwuUfplmm5aIck6KCqAlVRBKax/1OB6
tiRqtc/0+P44qsTUxVDOK5Zed3pGqUo/k1lqPiPF/51SeE2n6euLuGOWeZ2HO7BXvbbDOjDXz5mU
GU9ObACecaYwTpDMrJAFIdEXHPsm9AwG5yIHlm3muXoSoxXX9Is3h+qm8n56pMwsvmv2AJ2mshB4
14zJH2UAwSjA5QJjcOnlDTUpMXueGOpWzNtaVdxbN0XWVTIxsKuvKVeLrCwoKW+EskI6mNFtlyjE
JE9n/haIOnEOjjwExQxlab40OHKZWCgoW+RwDkHG8WAO7XA1SPOMLTSIfyfrVsSaeDwJiJ9FJB8D
G6f3r77OjKPPR0yOZUHNa6uKuCsaEJXHFQHcv4oVRy0WNTw3UKGveQoKh3t3sXzevE5l9rORM6sc
BiXFhHTNpqWPX5LXjv5cre0VpzfD4U0JHpO4oBq0iSOMuO39KKoJOuWSsvsNlu+leHHLooHD1XiG
2lunWb4dQcE1l2UqC/17EV4AWLezRglk2Ot7SHBX56H15iBYWxp6HHdXeeDtcvTJMS6vAXPZa/HF
0jgMEhVeiqtjkxPWjs4m+tazkJLu7h/A3xiuinM8biT77neuixY4QCgrvTLMxWOwfqIpdY/q1f6K
SlO9WHoiyxR49Q3hYFdhTL8WP00HH54uswlYYp7GqkDhAodbOfzke1E8ErAthLf0It3d4tJ8oop/
WbovvLN0UZPjctCdYocK54CAQ4ezdwq2fMpKEaAmzr85jHqa/Dzg2Bp1zodj76xNoI2qZSXXtkw9
SoFb7ZcLFb+Sqe7hViXxf9A3Wekhq2OwlYWQoafncoGGzm+FlqQ5ZvIUvwjiWlKYG86gqnwz5aBR
i2PPut5FSm5RmFUbUgJf+1SvsQ3I67eQoP04FaHzWiiL4F99/1O3XH9Sg0V2WT0pgADxatohNVb0
BIAP5EeYILz2Dfx3G80MkyPansvao/5Mxh6gkRfMGgrZWPHhnIy7JPaZaygZXpwcwT6yCO57FOR/
h1thSnTAAGQhhe4hXL+e5Mwog4MSRFjmELFa1w+phfcPLHJXwpAE1M4Syyt8yH7H3mIH5hPla6rR
zC4Xae9vScLwzGYI/u75xbmvydoCmHgSl2uz5cCiNrmB/GBQPIpByTPw8w1cdpyylAYFM2liRvFc
0+esjc97b2sF4TNbff78WzwINIB7reIIExyjjYNQZeSNjUfMeb9q4oKRVrmdZ/zzVTQppNv/ZDUT
tNuJjdfQeN+Uyuk2Iwwt/+IWKJQzIIMB6u2b3xTZRt1sgZQyvOti3D+0GORFJdl6Vean4KrYoI9n
uLAGeXMdGyjiUMjDsdvgA+qgWcBkOV77SfQ+1bDncj+LS6iMobD8EXZI3Y/ZtlRrV+Ddjf1k2I6y
ru/5JdhbBldx1lHpsF4U0/Jr5CptjcXmQTyZl30iTZrp7VlcYOvKLbR5MnlUK9xIn07tDJeW92Wr
CzyP8FDsDBIVK1pmBumhT0r3oljdOpAmz3s/WIydLiYvelP3YRzztfucZ5zb+f02xQr5N+i6Wxge
rBr3bSJzgjqJBb/T9jf6mK8hNCl7Vw4yGPN1eT4IEgWrUihLaYRt/+3/agNtBqJIKnzwdKoAYQbM
MG0Bn0mmx34xnVlJwk537a3bkjdMWdykPtPwpMi4M+1HxPKky3J4d/+miqihRjQqb1llcAf56mxY
7XlxV6ri1SCjoXvW3oxOnY7dOkJF1kpD0nHGIYUCC3UlaE9qeS3hArz90SuXMcc8/IfBJVzb0cWT
V70w79i54n0AFGtTLeAYWXRqAih/xwqq+ke/03joPBWoXNVaX36QhDHkbu3LlWinJCOtARU/jASE
v6baOeNAMIyUln3H7rkQz9cU+MWq3riS2Fj7kA1jKOhqyAWfZrLi9IU0JLnE8QjnbcH5ACpRsAB+
3F8WTmSGtwf4+kITFFvlCybilWDkEOzHY9RxYZdQduKK7R7AWSFe5fEBPyjmqRH+6LPBf3YIaTvF
Uguc7bIOtTwPqCGMnRTtKft9FPESUS6zTD/0bR/el0DXn3BD2GM8uhq+TnNPvSKmIDlwar1Lq7pT
7JjFDU2FEf5lp8NCOzfjivVLpV++lHDWlhRM9QXKq2nUNuB1J8+szG34XLAncfOmvMQJcPZNhpX9
LdlgKTr2hFcrOWxMDF4g46VbzM3ZKEm5glD+MZg0LbF0RFYQg8B514Kfa7+Ekvn3oOHjMSdeTY4W
eGWdWK5oeOgPeKZPnGE9tyEccNHl+wlsrAqM4m0pEfRXx0Y4k0RiSxswjaG74/PR4BxR7Sv19MKm
vth/XQXmXkESgrxkefAvNlEQ8bnzKswQlcqMLK5eU19Y4PcI2k0XsI0ua2U0htaxNGbSA4w40COJ
NhO3YBX/HzFCiT4HPxRM2XN09b1LQM78PC16APjfmovjCBWxlTMBgt2ZBecYecrGbpPvXtpxklzX
hMIbCGglad2tuUoDPeBRVRQthsRRdM+7BFkPRpd+0Tvip4xDcgKbIFkIppnQdB11FbhD4R2Kf8D1
+u6veO5nTqvcB4/yYKiTm8garr0ex8zvZebstoAWDIdav11FY/SiivWrOtzGh3ClgP8hcoThClXY
B8NFmsbqzL4G1Ha9Bv6NsyGVl+QoxvX3LPVOn43WxjLTX7rhAnvMM2YnqY8K8ruIY+6YGGtdk4HI
KTEtSeg9TEzmEYKeQNLNFpheyFSJWvq8P8FffkIZKf12wiXQZWwgDOi16qkxemn8KaWq1mPHgiYU
P9CE/LlVd0qK5eXejD1LB7AAkQJWDJGzrwYkLRHcLi4xzVAmX8BrdaKsgOTcBfkzIuYNCpMSV51S
hkkOnRHhi8YMvV/QUdhNSpaGRN92yO8BLhBv1apo3EIwb9dwOOsmIOMGvochet/5jevT+lDqohbI
EkAQhdQaAuVG6OORGxwqitf7B2nCsMyJEJWsb5B2q3EzQ+Y5R0Xy5jkcvjP8oxJm/l7XolH0NjJq
zFm6q62/3BnPZ/hNA83voa8XHQ2Yl+Kxfs+QIr3GrX4HaxrymSGjr/wrfZrU92uEEowtXYLyCL9Z
3h8riJCL8g3xYnhg+t48bL1OMYv3mVTeCerW2t0qqovfJrweNImSwRsH5XA+ucZLqHHwICUGMdeS
LUNIFgeiSM7bU/zf6Z5KSY8MGTYbtK2RSv5gReFKKSnAW/aw+0+REPzKAIXdRZE1TlGtw8A8qJNF
FbCwrSf6O+vc88tn+ZKeLpFI8ixvJChhrmCwF+cgnVbFzgrfFFVDlx1b9r2qkhD43dtnb/1dkar5
H5Qb0xDjZtUteRFZ/f9vO8sq83WY34STUF56eqOV/tssvFUdnLyj5cHYRNmrE80MJJGYkmmdJ/UG
PV0LR+c6XHrcYw9uLM/k53N+47m9gvir9gY3goJy7CpfKibfQsvrBHX78nU2a0DmUHlypMxle3gM
hvISX8mQBFbBwKobigcYmKF4ypaBF+BNRkdcJkabg45ABm0FMVNoCcGLLN6mleNnaEu5TZmtMVwa
cU1RqFA3cuLW6ssnmK3omJuMHtd/0E2NiOh/kcwoD73ceCEOUePpzWNNTpyMjYIRxXjw5/nCdJaI
vvr/MdwhMIwhWvVjQ2K0NjK1nxTTiTIZ+mITfPkQ+H6kq84Rx3HGXVLzaeBlfj1ONW/yeFiqcPP+
jZGpFpPKiCfCL3K19q7P8g8CIs7n79tXSMlE5e4GGIHMwmEvjq2N+r3d6hG5FZtZ5vOxhWV+aIdG
dnHlfRtxt4aqaYGUsge64rmVEq+/jzKkQoC6V8LM73LnkiTAbuCT3JayBWix0o8tk5hiKw2vKsFa
muF3GGNbPqqw7IYl67nlK3H6Y6GhDl2TSfZwvTe92aW3Om+30SWXrmmADbk2PRKHmPAKW40UX/Gr
a3f/+wJu6BRlnHcqTTfUIqxBDzCql4ipP804/K+kUkyraxVnbrAoib/1XtnP7BaqzS7vaP0JuXtY
zkk+zV/H3rUmTxIqUsVRMo/WeFdoPMaXgcQSMke7s/2KzbBYovPaLq66/Tp3uQ8P1mNqSBkr5eX/
QKR4gTK8cA50/QYe+/55bMa5k3MAe6NFi0JqPKKD5QF/uGGz0iDJYdBkLWivdPvNw/dGn26Bse2I
F/EDpSV9Rn3t/bRObl3xt2wEqdprYXqW2BGrXXvljrbZCnsj8yq/8FFizl0RIWDo0GdhD7JwpXqf
iX6TbySI0XmjZ/W3uOkLUHL4RATJjbBvxlKPQH1WXa89rcm5sDH1YbM9GoQEvyHZsmdx/w4kxuxN
RJGMoNsUSLmVwgmykSgXtPS7soBZ/IlObHWDSJhz0ZfUbN1BoBAHKqA5x4DyGTGII1d43bT7XoTi
U1T4HhDR1qvJXuFGnr6RFjdEsiOLLIfAB70WjuaGa6JP/sgshUTH7Opxze+4Tzz1ODxUPIMBHYir
OFQ/1aFnwVbICq09AGZEyBZT5M6T49i1ZmP3VBr1rxceHvV88D/8LxeUhyUKZL64Y6HTSxqFHpld
UdTvxmm+VE8hYGIyecIPKr3OUSAgKmgzDX1fc3HLzIW82rVRj5cpTpsPffQTmttQupCYwDQtqtfk
ygFaJZHYEvLQuanhH4uuV6lHDrGleZOnWtZzsdbDuVaTTdlL2ir161xF8NTKPLt+iS8pT0//Q+uq
f8DRGWuPFzdpET5tmOm3rrpNift/3Q6BCTPk6/gYRR971fd3auag3u+UV70j3LhPqpFkqGVJ/lHN
SwzenZIodBBPppEZWHqEbXgru3h7Er+TbtQVkqbVXW2j/qRu69Ei0LNw7xJXJAYk5Gywi+eEzwO7
nuWk0nR+4gs/P1q0LtpEq8FNZbM731ACYrNkY+bLbTZzg7EaZtyy2pPPUBQPc2x+ZuIbVW8NJBZE
v1lxYvJVkKnOCLAaqUs2hccCmQyDCRppUZaz1r/C1rYOG122KHmCKZ4SxvZBjVkA6QKJsy+MGNZe
N507nphg+Gj0e/MwuE5HmZ8YiEywGwQGyleKae8stLFTGDpSB9+c1oVwN3fh7zeBVtOi5ZUEtVH2
Zr3sqj0ePzxkEmlgdqZ5XBlSf7xmK/8aO7Y20hRVJ2KMJqWsa1SXSO3g0yxj//8MAfOfG3Cc5mut
RUZsvyAUiVYIvj7/9GHG1InNUxWABsZkInQIkJf2p0ERoLxFPdMTOmE7zL0rAp34kDt+egUQ3GA/
Xk0Gygles3KBb26byIYyEOcIZ3tvf8YRHY9LceWkpHhLZWD4dFPAeGbmivUc50s0HnShxq7OgRwo
7hKJ63F5LZQkV+F8TXWmRkxlyQlKeN52jIOhAnp9cE1Hu/ZuFnh7Y/lgXInOl6AxPWYw1JakyeSF
ZxCWWNO4wM2c27XXVZeypI5LyNwv/kr2iPYwtzid1bo15z/ROsR9LzSYY8npwtGb6fxg+J2sZN/3
xc3zSNPW/sNeNKCnJtxZ5ZiW+RotGAidOV7VMAJ8dXaBl6vJXcvUQIkZdsN2Xwxy/936Ftc5PkPZ
5sHJELaIKUq6IWNnWrJ42FRPqZAmP+z47cYulSiTCITYEVkI/GUCCmjOg9UJ8rRoy4yjVEEw0fHK
2XJgbcRgSPGjgSdj5CTn/v8VkfzoQSxWJmRzvMt5R3QHahVjjoez7uCNxHxDIDUleTGOPyLO+Aq3
Tk2Dok+zracS/jVrYl9SDkageR0gjbNseFtANBoPOgWh/c9v+pRdPngFUrfEk5X87DK3u8m6JxPr
6vt5wzJOw6jxZyABtYFktxvwPQCxz2WSqIDbTApR7jVECWX8Esa1YLTrWOhI8OlEEB+ALFm9aStH
fDwhwLO6PrGQpgl++rMsCE0oAM+hcyBUqmJrKq/w3mVRuvfiF5ITgCNqCcHqhcscLJoD6JUxQtxn
wbfMCcc39f4jY7l1/OBGi3ukavfQuOzqrl+ZknyEXD5ZdLzrNCLarSIzSuXdQZT6lo575QZy+kIl
rBAuPSB+7rAcm27kEddBWh8GGX87zQissk194SkvC0n2Ak/f4xBS6Md7/YyF1kbjb6zi7WppY49l
uRoFMl6Gv2qFm76Z5j8WdbZg2DqZK6+Tnzy70CZDqCzAdhKrsRfNxegg3uLX5OjjMvrDnfhPfOHW
NfzMD3mpjTP3A3wgpswD+pHFoskaXFnR1yaF5bhA8clZULRkdf911qek2BHZizw3CjPEcgTQNMN4
fzZb0xDiCX9PpPZ3qCAhiig1AaRDlnrGmu/lAViLhSbeT2JmoPxfZVUjvAvSOUAzERKbwc6JJz6r
EGauZZuuDP/SKwRsWOMrGekjivu4p7+Urt5es7qe5FqwDtYgf5aXlseqHVyKOr4zuAig8M0hfokL
TE4wQIAPwGMgEBn6PaesAp+V+qHyWk0SWMkXiK872x3sZ92dR9wBE8y7HcAKwc+zN4MhScA3VM7k
LhqGfXDUFuHhvY52TLlVJ8GQcBA6cbfqyQbDJ4nluKkSAJ9DzNxbvLcd1QfQaIeCeQcN8WxI9VVq
S/4jVz5x8TzV/dFpaOzTuujEUmZAjpMnZo+bLIX+mRlOjQQzJleyAbJIVek9QjTUcX6LZFZ7/eL6
A8OU7lSs/nWDNtJRTBJf8Qt1r75oCU44JLn+Ub8s4qTZbeZuo2p+iELsbdWgA050qPDFDFj+ePPx
xsfY0NpCOY4BhChOUTw1sGkNc7V3C2kiZyP+attA4M9HGh92gMpG+1Ks7UprSabqPPEpnq8HRtX8
BwpG+0DlzWV9f2ZBCbG6Oh40TebGRwxVBkmVxGvq19HaB2eMSZNrkdjYfa9GTftkb+qEr1J4DGKT
AZKdXAE0+h3UjLkfH9VRDAY1V1bbpxDsWoAS2NiiSu4YjzwlhrFwGVvVVYVehejtLllbBGHAR8hN
tb08mC1xUGB1t98NT/2atsAprC7C0DakWh9427xk8OWhUHrf/RWB5xa5Twu7h+8yzgQvDYAp3pd+
hja/6jcMxMO0CeWjVup9BP3fR0cewsYzmpduhFKYMPfZ5jrsx5i+V6eqq6UkrXPMiQbNb49/fc8U
tIa+L4GO7Wr/e1aKcqKiTnWLz9JO7+tcJn22zI/PaEmqbNJEs+8Okj9tEFSZV2TjZS7EWAkmGFHt
6PZZxO3RRDovqBBZYUxwJhbtklfko5f38tA6STBtg2HN+Aa3PZhws7jycTKfWWGOmciSIB5ejXqh
6Lip6RE15DkbhylQi2PyVVvT1TLfuFMixRlqm6KI/waahzakMHzTrv2bhw5XwDIJmoWwAtLMq8KB
0riOeF4MReGMQZZpd9xpye/KJLUDkRTwgWUjN3nH3iHpl/cSnatJ6wMc0AcIO819t79zQzBIHLiC
V3lfd9HHw/b7tG4rEaHjKNnYViiqvspDtMLBJt8axd5wf1vIyGD4l+tP8HkFRiSFxYpEEl3Oy9zv
Rs0q7tQUZPVtICrVbiNNNQgJKdF1dqqZ3H8wvCjQpif5Chsb/8049jdvSxI8ZIkmZ6Awp1xO3Gb3
DiVpAJtxuPhKOUCilzbPsdB77W5ZJAlqtE65LTKNkVbEqHgef7+0834YT0Lbs77LIvd309fU7i16
MfvFYVkNPMCo9INU/2oggN5hAV/OUr0Ukk+4lk+yClj6GiYM3KctUfyLbQY8HCIEJ8OOMrlollXj
RUb8ywsvHtjP537Ufr2kH73MTRwidpTtTIcuhwdZ0kcwB+K/aO6gl/4Y3Qox8vtIaMTaIyoHAV3b
H8tP3QA0/2Ovgqf7MTJdj9IjxvKQBpLWkDp/Ow0CVqGN4ZKefF/Oa25/Szyhl/dGqehBpfzmWjxi
4V/3lmFT2OXTZqgv6aUq07mEbpgc8kxNaeXETJkb+I995pIkUeH0lure/lOOMckI+Os2Mdfln8BZ
BrGiweYtykhiHNqxkw8OYInoWOKQRnK9YwgqUMX6dEESr3Gti0tMjr9SXxCs685kXmu9xnaeM/t4
POp9XBRgyy/EZFaMlRkc5UMlAfa2O1xBgjnHb0i1aL+IhSVu4Ia1ATKG3/ZOHxZTmY3vZkiHuqBq
mBUBUIyMVITdDGbqnW8N4zW2U6+jEZ3WR8BcP9LGthbCdBheFxXReB+iQEEoXok5baB5P3SV7k0n
3/tlFOYmZRSCG90ScCIQlnWi5n4GmVZYyPa960EN7h7mZ1tNFHZhJcafCpL8uCw0a9MSvDq+xZYZ
N2MfTp/3155G4uL/LZBPdt4Ftz7/M38J/yrGEMrBSOqBYj1WnecpiCUyzKHFvxmSO81Yob3I2Z2l
s8cvLUD4fjyMWrTNf5WB87zq8veVmY3GiUswVjcKEt6JgKGeiqliXfQugcAF2QRT2PmSKtc8Trov
Te+78ZSvZ16gC2ctMXOYstwSJ3SiDLyalVOPMtnYy2CKQJ8SWM68ZqYQ6m8FC+d6TQHU88MLvuVJ
RWsgV+zomriT2LD3ez6a5grZ5L293WIrE6klk92DalIPBs/ANNH0lZ2exHs60FUFsnauwljzffIE
DQ44zEhor90qJUaYEDzcfCTbXT4rvUIpKvv1+Szcp7TvsfGaIaNT689uPBbUKi7VOQKWM8Wcj16m
oui0qNqUErOZE8FD03Eeg8zPCfmPvETRnDnDosFepYZ4R7vSm+DfuK24vI9PUP5LKULtvWLPy7T7
lcKDCCfWJBI87IdkqI6qs+ecq1Hl/k1ew7iiCyMLRkjJ0ZmzsVV5zrH1au0XKtgYaS5kdHhqzIg+
9FEnBKSebsW4eo25i6gBzLBwETn8eiFwXMkSVRh3pLgFrBe30c7Mr6VwyYdXtuqr60uB8MqoqDvf
zcP91q6drxJeEz9uA4FDG5OoqzESjzsbR/Sk8X+VevmsKpTy+cP2A40Y9XT4nC3aRJxOOHuhEcVS
I48a+QIVRp3zLvFXcL7Gn75+2oLnhCPVkhUqTZOFZcf3MKIBvElHYBg4PUx/ICCr4NFpGQRpQ/8H
MzRZrZxFahmFve9wTc7J4xz51b/EFils1oEFfWu11fMkecSG1I9nkbkPBY1jO5S7neXB1YvvyG7k
sh6Elx3HchhzZPUCu8SrMU0UpyUHS9Rh8ZEu1SczGP/BZIvN7kw7XQ0vgcg71Bv4a3UOryEre9V+
OC7eQoqt5G15AxkRGxVkH5AdmGaa40ZRFlOvH1ZkYuCnPKlOlJWAt+DaBF3tCwPtaGahx1gw5lM8
9Y3Jd/toJnaKI6ApDnSGhyrXCCaXYwX/vBM8lJ63yBREVw7tNmMJtrjUd+7TqmdxblNs5cqxpSno
6LB3H3A28ZMX6wNznjlzxYrVmQhrMD2qRljfsWxjkO36WNMCpus2B2REZJbkmxfGeafWYqKQabj5
60SgPnXa76+zKzm7oa9MQvOGWohW7xaSa8ZL9LW6c0B2LLANODHH5OanMZ9s2DI1mHdY945ozbJm
zuu9yN40bIPVS6+lVUoGYX4qRQQ8zKiUYJoE2aDep9/p6xJett9OBMrO4/KvZL+trZ22bp3ZWTqj
a1wpHi0McK2PJWlpvI3EEDzFN605bi1Ipj1MxdL4a6iikJ5SNaRqqA1/+QUayUXChgwsUIzUgy/v
DPp9PzQXe86jQujdfLDBzfvrINuBHX+MyUPYafB+Cp5n5IRSpZfr39SEU83xrUauOr75ZpwCvR8w
Tp0GWlOyRC5u72NSDFF4v8C+dcI09BbjsPMdk2+2VxVc408wTEJA3HXbeg3kBF09jYLmxSYWG+Rt
iCG9YKv3L/9G7Y90wt/K8p9za6L7qwos76IkkhEVELssqAVa7Z5KEIWBGtr0sWyHTUJEZpCEqnnK
Vhq1VgerrE0W/ELnn/pNiNAKKZ/kuKrYRhiiIb/2BnDGrERuQK7yHju1ue14gCtZaGHg55drhlwq
BYgXTbtCTj480BswsZqolip0ac1aBW3tu7BbTMHa2y3RejKTWMXfMrCObmKaagfX9XXKv1pZazR2
dd2bRdLnRD8ZxL3NFXqwHIJQSJemtJ7gLFMSWrbE7C7eJ37oQ2x9WRozkXZMa0sLvTmWooYX78mK
ukoHMiaqA41gHBnVsiMQBqbLQcdjle/eCIY32sPS0YgMI8mlyYBnmOWC1ElqsB8w7vf7rM3mwdjj
0zAWRjaRIrD4/xgJdSha98E6Wfraus3ztm61QPA5Qt1u36/SGCgAXO/6OscQP/e/6o82bHXP2KAn
s7Va3IvV9VXZgw9yUwk/FwX0Em4Rp8yHlq2INjpNN1Xo4QsSnEc2k9/VmV1phTPy7dPBXsPkAk5Z
wLihhzRBh3EWxg6zLCEHndGnOTBCpjc0tucP52Ipi1++1T4VatF5/4+MACHWlQ+w32J2cKfQnfbe
bnXWitq/wGGEUh+OGftD5rB4vcG5m5jhV8ex+5qEzLXSvnQWmkXxcW+Z3aB9ehAQi7xOQv6oUryQ
HEXebkbvBRRPIzrgfG+F3M6hn8G3fVbKlalrd8/qDiPZMhR+qEvqfXGoHRcg7oDUmUXNOgiZUw8T
FMifH3/hWlayXZRi6GwTrembjWShgJ0rORgo5IhrdqXIAfD5FavbaOAumcDNChfis94JmcRv5cWc
bwcOa9aeOsESl810HGzKr2uOtvWJYlqQBt5Zmu9h+QAHo4fGFo+8cCLaS3UFEAep3xJAdq8fyMvC
qQl8Ms207qKZ00JavWj0MsOv3Ak4Se17YKtUF/Pu2hxn8QzZYhQuFK3mqXnmFYXdrz/0lCGWmxZl
VX43pj5avuy+mGPnpsai0j26o9EVUgjupyIXjxcn2OrvqUbXlPeLg2INcKoSa+pQtYx6y9+MMwGA
S+JET1TSTZcIvU/lcxJvNxKtkx3LcKZyDpdUm0JWXb8ROTNQB9a+zd/hOX7g0iUz+EkRLHjQ9lmM
Q6Yc7OZubRAlkNiuj6/1hd0b2qvKEZUd1zUDW4LAGkj4d6QAPuFdfsLVycX9K6aVm+ovUteMtbRE
CvtPXRliKBaZgargfXpvnDnwFDYsbVXDmpc+hWdkGRWP3hbNL3cOutMcNbgw75+7G7l+qRYtb7B0
EUEqlPckNX0KNNHvKOOixy1eX4l0cAQzeXi/hUa9D2AJwaOByr5MqEx+k841/IFs+E12CQXgvDci
jnvXkrx7ci1sFhvF55KmX0WE2wN1XkjIoY7RBHzKnmjgKSAa5NVN+FIlH/L1DxdvwjBHV+U3R5LB
bzCoNh0wq6xqbPysH1KGih/vDf54QcP/2GoEtCFVjS0rsz/Qrd1+jJiSKTuxIQoj4RCLzwjY82iw
ugLP+HKKwDD46qQnAelfdLU+PO3oFBNCHVC/3+4OljbnKfzxrFLh7HBW41ap5qabcj/5apIJcVm1
f2MaQFWN8aQRXehG1gg2fVl59hPu3wQTSX4X4/ujL/2LNvcOWNwTNWinpL2GXolfu2IS8Q8zXdcH
/XSzltkqpRxNu+Hj2haYNxNFn+jCsdg6hkoNJNnVhX5p/o+79D0d1NSNm5ul2ED5u9EpipwH8UdR
jTDVerRvEtj23+rFXhUjyrcbIT3NjkrDlc///oYkat+5tteE24Uj/1q3fquYyRryzQfRGIcuNe1N
1swaqJFJd3yW/0dkpCwHNwwtW1+mWJaLQSWgbN66V0BzIXUxpUmZ9TybJQpoDAgCTvu8eZqmk9sT
F7j6tJHm4732ngGCYmi5jIUbEGhJ/jzEDBUIdIp3TxLl4kWHRfmH5J0L576rMNVzt6o/zqYBsvAv
9vMwCskz3isTcbsSxS5io2e9AWPInb++gg/emL6t6aywM1V8g/He+Lf1K3KveKp/RRkpr6Q0w270
UxXkiEi3c2Ta1a0XnRQrjW1y5frsBzw6p4cTdxXcr2+VoK5wa9+UU05J1Qw+hOQ8vwo0T5jQKNUL
IA55Rx7dBac86efrLAlzh7UhruNhp/pcQlHI6RQTf/1vXm41QOByvd6YW5WrtU1iJfKI40h6cr9q
1Rm1YwaQkZd+umgazdBI6bGQyUuKzEjlQdDoS7SPWjSvISlf3pC/NTlNNRiq4Lyv9r0u3cE5fmn9
sI/iDtBuvYbc0axbzXdGYNL1AgRrKTKiohg5rnBi6C40SKPai4ZBjsmSAZTiodGFBLmUCcgLRKuo
6jfWlQ5xbHFXLdBSwkDxE+IKZFDunDZJ8g7ov1WBSDn47m5WlJS6qiS3mCUyLEuY1SZYAnyl/THY
Tn20P626PVTFm1B19I4DI/cJKBFSTonMoNeF9p755rF5Q/BuHi8R42RtNR/gW6jJLG8Vh3S01jId
Ckdv7oq5QtUBbWTuvY7JpBd4GEHvKn6vX5YTlwRZi4AZi7LYGiUExJWvMJIsHNXKVffefz+8KJ+t
tSUrPqnxExWCmiWYqO3/1GOaOJ5foPbISZh68L/gs35QV7OkhCVLebbDcjLzIGbr6G/JmenlCr3l
Rs3ZcmQTr2vrAPUXG51+VV86oBOQ5ZmuOeJASn414KATdJpajSrzTNyOm71mzYY8xPslKiwMRdmN
yUTRe9aoYYbi9ZSRWAwNA7VJYkCJSN1IB3yTcXpiNIOm8V10pKzG48EC47+v2V94gqLVzdWYiDw4
ANFerpqewpgf0y9oTuAYuI5bygjp0DQ+3HJyW+5P8YpKLmk53Y7loopapoHA3gMNUYntSKYHVWvp
W5vWcncUb3oYsJIuHwFWkHFtY7zRix/PpW/l5OieGl/teD7+VQi7KUeVaEjWWxUg7jBrDlOfwzaJ
WDpchiBlhwfc3ku6l1fYD/o9+RmJsjzVJxZeFv5BIm/IzdFFX75htSvHfBgfIs7MpqoZcRuHKlsp
brk5VtBAAiFyHt1McXkVaVpbpTT7LtbIe0klEjuP17tECJUpZ8cjIKXnH2xmNkaCZGziIH7NQMln
g9XdjsRgeiD4t7+Qf7oScEahIIJsZHXlka1mHtKq77bTcPKfI6j1TP1tJAtV0ac6AEzVE3azbRB1
S8qVNBU5zYduRgZeDmqAWK2WT60+2GcG+ZHNYgfhQ5Om6HH2Jki1COR8N3K+1IQklMZ1QnSAoSho
pmVS9IS4Lg9CHJuAsdrPfdxIkE1Kd6wUocYQ/pgAA1YaPwN99B4bPFFcHAcuUAj0iZdzfRe6NyGR
UC92oQeMczDC8WnfkS9QvcgqzHKJzCORXdpP6zOy/2m5/n5dMSuFK+snyjJ7IvHroq0UIHbIu1qp
Zv8rfk40u7a7cul8fALE8YXPF2dNu3RQ7BqELV7JF4jW1Lp/HLOGMR8N0kcAyIAdFoj1HRzmY95+
iaE7USiKYfJOI/qmZAyMJSjtLeYPcDKhh4MRXL9dk3OpY0QdI4SYGt7Ii3rTJM5leDSR3U4dkcpA
MNwRZAeSq0LnYejtUfVatzBsDPM5ldBoqBIE6pFXkr5AfPBEeANhWbyysZ7xmiiF3KSi9XnM1OUg
umVQcs5U8EkpAf1EQNxJXt0AC/KJhlMuPmKt4HAwpMsDOSuOhYN3GQqrIhHKOtO2lCPqi0CMB3ty
cpq0eSUU+mcNo4uD/3rednjm/cKrmOQCvj3Z3UM3hWmKZLRIjngJEbpuxIQxMWVSyHqMuCoWN729
lxHElpgVuVEH7QNJBzEKPMp9QmU5zQbEbsiQM7rQmhZrSWX/qUJCGHDPr0wFzSGEUDG2Y0dGYtU6
2gCPqcQi75MBvIavA78kVfHEMi6NIEiITzSxvJrjjxXYV3d3EjLoHL/N/rbjDmEWyX/whZuo9X+t
oMKUqN//K5oFPXj997ELkkZSP75B86u9mMvHXrq4tt3S+lMcVfdlyc1T0ZKVHDKmnZKGSMV7X1zL
x2P3P7JTdq8F/NGYqIMvKQNXOEtzj/aQIMfxsHxpHPSop3FsCNktGDXTYvestKhCkYdgaVeiCYim
4QQ182JVblj7MYGf8MTHrLXM7XVXJrtiYPXzq3iS0BktyScUfxPaWJEtnntgHiryTujEGj15pRE9
YOXP/GynCOpnMoMUjUNWhXlIaWV4xoEDGZkJli7oZtav6ZXA/e97PKrepHopaPz/0dPfIdHxwzQf
qDyrjNZYHR+WuHlCULhRV/uS8GmWjVQB2RnareB2U6g1l3+9FZUACYQefxxgVEUtWV/dxoF1hZGo
prNpjqcZ/ej6CGFN7z1eqxhi0CBZs/NzVjBnIo0mL5kQuLwq0clRhvb5lcgup9xwHE0CamtRfd4Z
xSZRXkOhjL/QPkBtTnufE0+upWHo3Y3DY+GShwHkvIM6Xg+25kpTivqQFoCIZgN521Rufi2Hf5B7
dwu/vl99aWAOfAFrpRNds6jMuQ2hAPjAgDvtj95/8NFfEkoxGONEQ/gpC1ZtytbnnwodeFYKnpKx
wUgNtZnPAxkw5S64ksXeup4338HN+iLOTovzVOo7p4wHXqGGGz6pIji4VWF8CaP4ZjWGS+dHn3vB
Q4S/ujjFuWmkx5pEiKAgwXKxcgPeXJ9e23mdRbAAY7ZxnlU77D9LHUZhnQMzB+kCLVP8YdMjziHm
EVG7LuZnzrnu600CkpV0amYIcJ+GMQT3dk4tJp7hP2poFG0wcwqGjPCULuAAZOF6NzqAV6UC+PrA
kkvXl0Si2g4t8Qc9GlpUcRG1PxGqMfWwEAJSyOo1e+Zjb852/HeqVzHdZBTT7SGzJq0DZoRytBk+
S2dUdfaNdKoKVxcOLMZMb96LLjH7OFSqkRtj8UDZAgkUp459QfJusLJXbTW7WUHnOdAO827lsyz/
EwQIf8nfnxnPnC1IjMMyGBD6M7RGRuKboHBMPOs092vfvcdF3ENZP+PbTYZweNXcJzxGUbwzMYD8
VrxmO4bEJJgjEVqxqurwxc0LuRDy48vaVptD+wjxllwREDr7gy5fN9L63lb2EWwGW5OcOvoMsPWJ
5+OLfjlix6R1yOnusyvXFBAFyPZCubVvdyastxKs2FTZmqnfkt7te0onJeCsNRUsfR7vEHh34HEo
9gr9tGxm8F5UNLKgmv1nm+3ZkO//BAxtlm7ECXj61J6L8WoOvRMqWNPzInX5viFdUypIUv9ThTAJ
aPrBrgBb1mazt3E0SY9zzE5thh5EcAjUvMHnAEZ+aS5AUN0PpbKDdpA92rBQTimUVB/QC3nZl2cI
4B9s4WjJZH2H9GIvA1VB2+a5+wDTUaWG3SfAqyapcOwrRNDA3EWfqz5GuEhA1+VFWXCkdeh8+iIq
7U7LENAFgfWTGgx+omQs6M1LiqSZ4r7vMbx68rWRsdajcOrCDv5P0+7aFTaJcGIA+GV2t24YBMu2
ttJreydkNsM0RxIZBWfnnZnCV1JxePX3zqgvUsv7UePV+H/7USMEDAltD9hdBEQF5cT7hKNeugny
A4mGCRUAc4iKAG8/v+dqeXTWd5KeACSKIg1l+hoXGqnezzE90gffJv4Ua3lQmUrLtUfEyssZe4kG
+C+AYSowXpzQv+WAFDxvJOxHebqC/SJg1lEtIK3uFkP+iVrFC4NvythDY37pPaVdJwYhDcPxZR6p
fylnioX3FN4PZ39wtwu1shI2cffQ11u1do5OrKqXf5+q8hscfp0Nb4cbA66RlaQvX0pAeGbS76dc
OgymkVULZbp5/bf8Z0e8Lkdyz2jsc2/+PSfWqQEiTdZMaAIii2g43bwtt22I9eIWat36R3hMWmP6
qrdPicQXwjXtdFLXEuWh0d9OMSgE7GB2T0eOeeAilazsnsPHP4aD/spX5AjAHOCz5CQBH8NxDA0e
vMvI1YngQQdHTw1pmHlKNqr8zHh2nWy0IF2UWG+d7PHH4eonjmOJ43EN/kHU3H4Acy45HFkaolFQ
1J8JjVYa9HcgYb2eoB551Q9CvtLptL/RbIm41yTH0OnS1C0xrrten05CzmgkFAS7IHocdbG+nUtv
q9gwCmUx5zSgjrU3XcQmnl6Lbz5gSOY8ePDEssShbROMNDBSJamXk1K0fp/tIdMeQBvTEFbIv7dG
qPXVfjJpE5YegAV+1U7fo6dyG0HuON0XEIUMYpfE8QeKczpEw3JLpCJdM6dHwgbZt8MhIWB6yD6Y
RtqbdtSIV3cnZfD60b3qqhEEv+99EPxtEELgB1FaWmGkyaZ/j4dvGj1Pc7gnKtkln5m/rFpHNpCV
x19Kx0uEsiGQ+UVXiEQE8cQE43ABW0A2tELrXj9II2WFFdSZtuU5c2Qpw6eLSmZtlqzfNs5AFKb8
Ld+tw7+hI1USozeztFSZa/copEe30lJQR/DKq8XmY7juXMdmvTtfXzdRhuSKXkQDmtwxyr7ibv34
Y9dBCX21lh8+mP/+bjW0gvzzSXHo1R5U2RMAwaJXsWDxn6dUkl0WdLfhTQNgiqHGRJsnaRgzONac
85QcAoSiEWSm9pyNiJaHEViy/szf6zVdFt5PRAeVCJ0cSvIhUTmYT3/MMmBZ2kj5DC6ugvd1rvNb
PYOqakSZWa5B0jOZIsGOw7rEOnuk2Ex37hZmHcvD6Zun6WO4Prq/OPic3+p886hAK5YOEWhqUhOj
qHpQsPkVhkyFVKjTWckoD2ipNYpBEADCK3YE328PR55vZp1VWAhVV/WDKX0p8HS/T0ppcLM6URMr
2ONzHLWLioIOE2M4J7UhhApB9hj5RNU4H1mvR6Yu3ZwE63Mcn4LLZWDJE1nSsjmd5PDBiBE+RdqW
zedEnH249RjeDmGv9e3zIWiTQarvq3TKiGj6E6R9NAF9aOb9++r2ncv/6W4fev6uICrcqvtxfKMK
dDYhNSZiJtKDnIY4tsPwI7q+hrS3JWrpjO5wr0cSEdOnyOWECLSdi5XigE27GLC+0oZtgftYD37h
D8lR9SPRtm96gCjEWljTF7KnSQ/PxbZK3NvrMp06/S2bOYA4+jNAoBxHksG5IV5X9UgUlSh4d2s1
Xg7HDyEO/dz+8sgjG124i9uEw5cYeuzwaTKclky8izPtSM1GOFp7hgIGEhznvGOG0ntsSPX6yPly
eX3DnexcKQeE7SJKQWoWlspfN+IsDxXItkVV7Ty92cjnfkZrnvYnM6pBWkgPQ6uncpXjI8GpSCjK
RkAlwUB6maXO00d2fn3Cdp0t6QA3AgKO4UkUeAvMdxuXYlGLn0yeqMaMKeqF9aB0ZEWwXCocxyFR
iF2GhLA6o+fWqvgxiv0mTAuW/EJopZhJFL/A6mEM4nJkDkHsSqNusHefkvku/6ChfbaS6tKkUBZd
E3AIkdk6tV0VKyj7eQKa6KRK04rNJBramWw73IXzmsMSKYES9Ch/oMPn5N0AHsJgA5H7S6II6mCK
VC0M3HO59DMXCpFESE+/d5SVrU9K0UwbXwn3w0niRiIYZqyc5wA8sX36KEGAzv2RwnS9yhBpa1sa
7XuOBq+Ac1+Xh0GIr4vLq4TSrcvyH4AQigoUeLef2T91U5UAZG7jxnu1dqp0Ew83u8piDOj3ZEyt
8D92Gx16vNEWRqW3IYdC3xkHfvnJyDwFhtR7iZXi4xhFQ5HCS1IGB2Nj8GhLuOkWRr/p+kG9kfGC
E0xr6qSC4Hy7E8I0Hk37GbP/l6RYuOb2d9COesMfc/KVFVHjqFKqcwOwZQJaSEXELZp5n9q9Quza
MtB/3Wiw9xVs+hy+a3vEQ4Vg6BZbA5IUJuNVdI0EOzZg0jGqk2srV2s++HYmKvDNUcj7kAbR3Jtf
yXzDCQUDotEOX8ILU3c643BptcSXsvwhC32IVPBzBzCQeUU/a8DWliWre6gKtlqLTXtvYUc84EtW
dMU4KsEp/F/N7m+pg1K+390K9iJ8iBE5OjvNxidihR9neHpY6hzl8w8Kk/6U1N/+3uplP502ZtDM
R2q7IucVRf0Y0HH69/TSHCBNGb3vLYBCtowYxONRoL3oluRdjafOhAyGLRuuGDoZt80JfwL5y/cJ
fWemzBFJ11kV+zuZySoB8hsTzxaSNODDzwxZTrNFjsX0vu3I8GDwXTG6hsa+rCDuXJFCXrJO8yc6
dJQONfYP3EPzyJuTVNafgPZv+LWG1fPvLILSNZ+zYnMEImSBbkX4UPgb8uvjhgRSAOXJRpn8XNel
gojCeNrr32PPWS5Z7rW7nkvpxIsSQJsvaHSvwIo8y7TSATJ1/o4MxP1vnQDiLSay3KcICYECkZwV
0pALuYTPHlw+oGBbr6xXE9QS+a4So8PlrOFB6YKnFK2YSB0USeol8yLBI9nkRu7PixpjpCE5KSiV
8i7kUmRO+mfsoOZG9ua0/NnlFWbk1mrWCWIc8ANyzXf7jf0HY6bAkYxtaDES/Ixo9FLbt1oBXxFd
vG2WFPBsOeGnz4WhkiLaIDeRh5crmOn4iTVVSt3oSg7TsGaehntMkijRAuzJRpkWonX4+osRn5JX
rjXAWg3ZKcQBP47EExHTc45MPqi6yhAzpMACEyZcQGZXFY/zFmO2Uma9BFUIUNnRHoFpbAjAvUal
IkjqdXPI0E6eit2Fu+pPra0gNN9+UQu7RIteAL7SdmDKRKbs+X9trQcARqVjwPvhRYp2JMsgfPJN
i8FaWor8tqXB6VuvPiw4tMZT/DSlpG3XE/V8ZWhIXzxmNh/rDKv0uIsUDnGDn6EVWWy0DDTB5thu
9GdXK7fQ6aoNvZis25QUYCgyGxEMXR5h2rioXv3I+Ckbyrqoa7DRR4oqTp+rCehgM8rQwLOZVhzb
TK2xxswBgJNxcUWqBqLYowJJkEIpgsU+cXJ2ojNRhYR6ziSJ2kcdOV2ygrwHO8qNgZE3Nk9PyGHq
g6WJ2rqD5fHUVA+LezA0YCfl7CnzjZLgjNd3zMYd3thRRJ6P2PqCsCwxR1xFR+ZrG9C3UquXKV11
OCwPbhFqaQME3HrfmZpMCWBghOgoE0nA8MNcCYLSKEmNmf2f07DIlzTvUeYWjVSlHTgDA/7kVKVz
uJdxrshTCPudK+yK/Mb0Ge/7UeXpGZpmvdKC5fZ1UDpW22VUNH2UV79Zg8MV5REBkOVa7HXKX9yY
WYb4En+FDtHVe9uzyywVceadkLF6RakOEFCzsxs2GAfcUZCxSqFKdNTIfBCd/U6CBqVUo0VmQayW
BmQ1nEshg/k8eb8Jr5oFYHJbyRVUZbtbrmP1fMhLIcAIpRfesupIZaV5CMgMf0/yZpmuH1+p0FRB
S/2nvM0NWRU9BE2RHjJy0jgtFk3echUl6/PQweoXGEloti59EMOecp4e+ajw9q/6TA9nQFb+CwBA
9i2smJ1BfrV8+3hHLBmWH6+q+WntQ6sZmu5UpMkoj5lfDmpA1QWcn9x20ltCXOUuLGSGWqNysJVN
ENCi7dNuvfWeVs0fKpL3aokIOqQZ5fYtF0f3Rk+pwbcwWo2dI9tcAjSZrUzHt0F0y1ip8lfSb2fn
wD2ZkNWptfc7fDiE3qTWwZKputETBL+nWkpq97T0tftaD95SrtcRy6NydPQZc1bKFs/BTXqcU+Ww
/QbA593OOs3G4VDZ8UnLAipNjpJmg76NsCcF+uAA4A1TwBPqPyjlz+00lxNq6e+AGfP5GL88xVrZ
8MbnFLLDEtZRznf2pcyJEE+Zo4UtXlAAEg7CTurmQXiksWja67lqWbdzBtCO+b1MFDkRgCTt24Ad
iMnNPKzAIF4Bkm45gV5qUy+3fRgCXNhUxoiz9DqgNIRb/yonf1mK/S4Do9aFJf9SeSLA0m1w7emT
3BtLCPU1RtE2DpP0KXTOTIUyKw/K6yPjdWQLLpi3qMIw/KwI+k3ycnyk/sDQKdDG/4Y5x0P1TM2q
rHCiBpaJYyRnQIk2MTBy+eAnTqFKO98+CFMXufpXXJjvTyWlUj7bJunX1ALLpyMwfKFfZJhqhPyD
um/3nOz49s15BK0b6TLEGmD7qcOG4eNGrxblGlZo6qwlkz5Bj1S/siDsU0beSxmlm94iHG6911W6
/cnMmCokBamyLyCa/9dkxZ1rjHeieq3npIgq1iqbLrfDVyTYL596KCCt4sfPLAdTQBsRNsVmmnJj
tRpYqBnzb1G3vn1/1zUveVHzCFGtusFU1UBg/CiivyXKY1kD3fqcgnKn7Z2WV1wgoIeI9Zy2mHFa
7MpX5kGAIehaty21IMUV9b5knNfxu0S3sxUjtgYonU7zbLFYgpaA6cOWHJZggnyFwwVA45KHyDzJ
fgGe3L/dqdbJdpQ8wUNI78ZsifMzesG1YaAP1uKjFkPc+lzzbV5UnUMOX61ds55Vrvdu2yOHkp+X
NVn0SPoERydbmHaXLiccOD5uk0Fa5b/icwsSopnnbYOI+HU1X8Cs+4X90+BhLbwanRkBNZkNefGO
cuJ3GOEEWXjZQzd5NzjI14XNJgGX3+Ken169YLSV26iiOhW/mDp8ohQuMCVyqMpUPkUd53N3Bv3R
W6u8YXfGPpgCPn82WAzrpd/Ca1LVinMQSUrrcipNk4IluzDULy9+9KlOu7S4ZSrdOrkGnc1aq4KM
FFbB9YTHC5oVglXjQ7Bs977+1vxoiAnk9FCEY1pEWDu2pTmTXEs9fMJTg5eqecOZiDprHvj8BHDG
8NdF0vPfH/hsHOogHrO0NrrhwJCR0Xok8UBGJINUGm6dNf29OBvMNnX7BNOuL8HM7rrb6aaAA0F5
oTI1GiMy7y24bhWqLMm0Qsa9dhNWojq0bwhtCExPRZaliGNImMfFo1T/2Zm64JRgr84K7wh+kCPH
vWe0dgF+92eYx6NzSw8UK3EyAeY41/cA3ejSiFie0lII3upEnfiTQAvdCoviIcJt//My9GdWhRHA
8AcPi9n92syQsdFnADOW1yImOQbAkcUL4bv5E2sbDdYfnpy7sEfGgdk44nq5ACnvMaE07a5Mp+rJ
yNkeWFs6yQaukD/g/VlPSvUX9fFYv7ja8wVtj07PAOp/HaqtIbfKGrDeG1FahWyPO2diwgTUobZw
JvZifLljbLGbtIHf5QTwj25xl2UjyRb8Keggdp0wdfE9ORJmOR/NcXCktWeMe3BV27xEyRLNbgJa
uj0VlzgRyu+WSjVv4tcr7b7Bdt9DGPgcqFaQXI+FqUAMCFDdlTZIhGZb+hKAXjGpOZksVPrcSVhS
CyW2Qps9An3V3lE/X7nA86lsQUFW0ldyR4+rcFSwSFqwVEd8l7uLf0ThvGo/bWsAla3acOoy+jZJ
jUhB3XPiWlLzj1ZTsJXGID5oTRxjftm/pmHU7Euv9EznVNY74Ecr9z/P5qlalIO4izqKbG1+ZU/w
Meuv/KLPzImRywB7x/fcFXnIQdxb+MmjUdqT/8Vw6xt4MkZlaxatQpu0IV37wtpzokBxs5KvZeIk
r5ZRO44domkCMv8r1X9CZlOxkxrQQQEsz5sLGPAK6dQQPGdUOS894LZM5TfpqhMC4EP+AZ3l4kIn
wSOppFWEAK6RKiAKyvQfnc1SVVSPR0oTiwUaBlxOJm16FnJnGkx09EvTS7UxJKrKDLdtZqm4oGmP
oNdUXTZoIHigeJnJBffWHXAgdADJnJu0HvyAGMxqnO8MfzaE/8gCHvn/+0DLgEEBd7UaFIR0XysN
0tlu8K/S0kroxLI8EYpk6LZL6zNXNgLCEgV916R7uX0MzUtLOKVMOxQ42S6AyxvkWRbFNkO+Rz8S
S4EaaokLd/GGIksHIWgO9rLHORYXdCK5DZHtkwGNTClSyFV7dH+TVZNxt4zC85glEKm73PaeZdd/
gpCLo+7CbHXkbJBAOKn2BQCK/zMAZ1EAyUTi7JNxfbvNCc4qaLR7qB2XDG2OImtEFUzUnkANUASX
KqNISh9rP/7+bogREeghQw1ixL3MlExT18Bfyky43hE2u5Y66Trjq+hXYMeGy8mYfxiDtrQd0hye
Uo7kF2ZszYjhTImatHD1Ucq2gh4bjYcW0k6sUzucVLu1eBWSPAhQHXjZOayWTqYNhmcSuwBwEA9q
jJXPEBK9fFnF7/zYrWNk7I0kKwPlgM/n9OyGKJ6ulKlY+pQ1yqacMASA1hCMKiV0Oe1x95oUW4TX
uD0nKKPqg3i7WShg6C01nbuuy2pvXlN+6K4qkBygvJYx7IRWUxJuKcwfmgGUXnDHYri5jXvBsJhl
YWAC+s3pYTXxj+f+rmsaRf5iBGn7122tYZWaxiIHo7dNsHouKgB2pYfzKlv2s5ARUsfHzobeYBBD
4v74r0mEc/Tccu7L1OQKrE+KNYO8Oxnw7lIyExeu36iB1xTAx9RX//RQhDeUgkBiT2j3lEWAt5+M
FhwnILGWGCB5D3im3h4pjImnBf/DFLikkWqsp2q8WVXOxMhxc0fYEuEqx00Oqd8/CuNnJteWDIwN
v5AchI5sbc/BAIAulh7FGKFZioViATck4/jzmqytUkYYv9UGXQi/qY4PAMWn8cieB9V/4oTmgVL4
jFTNNZ8KUl7hHKCpN68XdVayXSPBCcPYI/8bZs5AQ7Qjn5J99ok8udPvzdZ+Rv7ZmtnPkbYsFc2N
A0xAP8C/AyRLED2VKoxZSHuwmKQjP6rSXL7a8JR6nevFrfAu+lBMjvbvWM9DdJJGKXr+ybQutTkL
ueTKvio2+jXAFssmNFx5djPZqmwE6+/ew/JXEP5/ngziV68MxN07F8+vID3+WrbJRZfil0JD8o2m
P1ExSOfslixff6uuUIYv8AGzS4yANddbc26UaMNX+co3TkTUcF1uWhVtFJrFbSB7c/UQPc9vv9iA
94SznfLHDfCAgQmOex6lGkOLG9UUeIrJ+x3zxcAXbJvd52XGvOndtru7VsFxz+3sjByOcfFcT/J+
PQ7hX3Yf3X5i/7kjqMqQEMJ8FKfo5HuRPVEsPshJw8evTiPYad7MMOclQaA4rK/mVQvlPLQp82Lc
VYWMhb8sNc7xNEZMO9DtEGEYY90LOzurhTbQTR2/k1bI6vQmYIf3gmGWhOy5z7SHmgg4J5Se+Uqe
4nEj5Se4m48BawYYeHi4CFMzso0njBE+xEtt7GsARa0Gweex46DuBNIqqY4GQmxmd7V+0OQnXYue
dj9dxp19ELR0p7eRySQckINxQGVyQLQsphlr20Ecq4MqtbAnDWySXw/WHbhHEd0cX2fP85H+H5ew
ufWFXakMpsmmkB8WWEwDXW6ycT3dpwVC5N2DINY6a1E8NVIKROzobANGIf1usH8sKMSjWCX/XJrs
YVosMg30TpjNFNIw/VrCKc3QSPab2/2DEIlasYeLY0aVMsVrIuW7IHxI3Ki/1PaIyuiy7r7RIwew
IiN3KFg81sG/Lm/cT8J2Fs4xWLGU6n6AlLGZ6O/HZLV+yqJviTdm+m7hNo9DkecsdI9qo4YSC28S
dm6H/6W532juX7xSCXiNyQTzdrojI0F/7u4caNqTJI5UDGLdeoHHnz2m8zbRsnBdPgs61Dx9rxAt
DQxUG3amXEWi3//df7EIe8tsSuL2AkBAHMBFvJxJKgJbOYvDJ+nSCp+V+qhLml7+5F5OSABYG6Tq
UUVD+1mcQpmtZfwjIgIQOsaQ1UMo2W37K6WpO+E9gEwpxM0e2oEO4sb50j/2PmtC0W/Y2GS+RnNa
sCJfCxzZiU9PR4SfEEKklRD1KFV3irVfth/JeagtNHCREXlHw8INleJMJ8htJm5st6923IExJgpz
6Zb81JYI6DNMCnsxvVAe3w15mhJlPjQTEk+AAsNIH+h3rRPF5r1msqO753zoGST2QrK+f7DodQQp
LWgoIHtT3HUW1a73RjMDVjRBrz9NneRiYsHkU3stkVpbmq+blUrNQxQCGc4Fk/toQZIxOaiw31oE
tBeh7m3EQ40Zuv/67BZXA/gbILRaMzfVToCU6tFLMWvWkxYE095owfPggtzqsp5hM5pWxu8Ua1AG
SqSZ/hKR14mdyo5s4NHYO1DIu1v1GsYLq43pgEJFaysKjGu7FGNAdpblmJn08Wx+mH8YPIf5N2II
o0WquMaUi5vshXE40NU7J1Sx8JZDIMFy4lNimiI9xbeqSZUefca1TpFYmMGTO3VNItxc2a5vOsJb
vvTofsb/Bu1qwFN1tnQxmsLKN07+uNHPhWNWbU608QI1cLWxgKnG4ohSbsRZoaobeJad31WGhECV
oe0/vMh4VNPQruKXillkrL9BlJMhekadeN5Bb88mpiX1dJ61cem+YYXq90REmbNkmF/GixxoPYF2
Ly0NEz/O2gqCV0auiq9JFxqGs4N51oOycPQS6nyq7ElwDzNYklirt3yF0XOvzFt1E13vs4XBTdXu
7M4HhB7bMpLvIKXfNAx0cvk4mBmGff86rD0Co68k5xadJSN8eQmzmW8msZy0NMqzW6LD1Evekfw1
YwcgsZcZgBaYhUDMto01hScJXe7bNk85J0LsSROhnnYNJBUAyWWyant/sXabpkFa0w893f6AZb/r
eT/VWZuUn9KjY8ryaF6b4V6kvRvd8f5shv3tDiDvINtk2G0vFmgfbq/Zl4TkVkxl1G4310s7jNUw
7DNU7vyj8C9KfsGA/B+S9WtTwefjNzQtXhwxcRo4mjwITR2+GlrJccQhVmy3yXTTbkzRbFgmclEf
MA8D2SOlDg/7z+3mdpx3klRiKrobSmQZspBL7n1H9/XSr6GR7/wjJWhVVXGxPNU0KK4RY4KcvX5G
WkPycYdYdJqa2p12dki/F1PMDp86XbGCWB/oD0dPc8RtGHtNc8pReZt8PM+IludJfj/sVlE1e2k0
1BEbySti8WezkfKfROB8k8wOiqe5rVJWtobl4cAhL6eXCMkWsAoeGvZUKELlgREjA8i7y0WNvUXu
XXxjZ/e9U0L2cJE2mcIaLedSzZkEtF53EiySbqLAb4mFOELhS6qnQWINkOlLws0SxE+2Ga2LZ92P
xUq2XZ1kJmR9o5aMZXNcZdl8xAXQzH3DoOpOUY0ATZKVeuJpAG8nCsR9b5s9tq/ST1U2ZxKYt5rS
LjBkzVsAsIb2CEm644rTUGAcMJ7kc0h0SQzMGOudDH5W8vFYk/vggOiYi4v/tL1IbMSnBCaM5Pf9
CuiZXdTOTTiG4+y77KTJjXnaWiGKRhDjQSORQf9H1a3BzmOVq988z/s9JCotFO+lZv5UeQ5+n2mD
mromipowQs5IdPdPT+Z1fgvJBfbrVJaieeKhJ5U+L64Gx+W2eP2Nq/qy5tc8oRuWwD6eJ9oYh4ZH
0w7IoOSBlnzCZOU8v7WIKhEZIGra/bdsWtODNrErwcMJ7JqENs1Hv59aHYfMoPSariwOeVyH+uTe
NBkG5lBul6uvgNnb00oUR2hc/oZFfE5jmUWZlzbtFUQG7p4LPjHv2jyB5x/0nkgUeHsH8HU853+A
oVZFXwmVSldmFs+5BofMI8T/YFkbUPnH/CXmgp9rMgswEq2lBYE9s9MI6zWE4K/3VmTQGHdzqnVZ
Hz7GdZDP4SsfLvahO0lnKBDKa73aErFodyIMgjNeLjtebOAxpQYXEZtKSpw5Zd/K6LYvP24LWsTl
lUOxiqKg1lCZM6zMp4GMEGAgb1dD68FhXMflzBWCudMEJXdJuC5mUWxICXFPLPyNJGdSy8DHm2Mb
96+Llcwvi8Z8PZO5w3Fzg6enEGRniqhbEFrwBTWeSg5FJmN9zK5ksS1rmGmWRF7yxqzkDMpJ9qkK
vadDyynrwa73XeQ8SbM2eJMk9j5bwftfb22RzTd2oYlCcGuIgDb09O4UYzCDEN0RFfBjpZaZWP60
0gHu72ljRO7CAwDN6uTnSz1fukoFZanFDBNtmUUGIlFNeQ6uGj5ZKf1Ijoc+dFhO3Y4SMBeHXbuH
e3PRCn8Nfo7Xz8kcWvl/2DJJwdyafD8yz2h8yskwdTz7M7xvys6SvYrQGr+BAUQSG9pRwEE22D62
uuDX+qW5J4073Q4eMndb3hc6bcoz3wOkxLzsLHAtLjjYQeI5JQ0kYMhmbeBlIVYX+FpWqvgkdgLQ
aNhQUtEI704Ctxl0r7mIPObOZDtWsKhWdupHozWJbb20v/UMO6Ju4lPooFaJvoimRPfZWf6WRBcF
QeDp86r+iuDg2VFRPS01jk/R1L/pOHl0sekualzMCXy2hecarBEpS3skwWvbkHpMsMtwQEjfySNn
+m9ZJoI5jPkuHvwADC2lGmKoaaKYnGLFMRDct0Dvdmn/zPl8ZJ3snHG0Jdkk/wUmURXmjPFokmff
wFgNGaJ1HNKKfzQBGE9sgvfEtACZ7puHsrcNU3WqMZLSXyfuitKDVxfH3rlFqNLmu75IetoUoCsL
keYX7ir7In1UnXg4NTYCxfCN2MbL/M9UHUKYdQ16mWU0Z8cOTi8Vs87OVrHRUyvbiEzgi2bvOLrN
h50BWGzkSSv4FU9YFqZhsFzcQIQeQ5LUR9D16Cmp/4ZQe9SamA3lwkZY5QrcY/DTU2Y7H/UskTtI
KOKaZycQaa+pPXyYsFA2VhN39zBBzkhD+KpcbI/IPSP4cS0pZJvbT5SXX/OxQt7/2VbFj7DvX6GT
Y374o/yrUhbCk6q8eDx2w0YLCb8yIhhHUWBfkYLGxEhSu7XhImrNGTobu83UKVBdeLd2j+5/1srV
kt0rxR+Qd+FZYLOSwKtEoOWiq9g56JjSyvfr/9CrkWTXd/JxVSKuSchCJkcO55dUPS/0k8zecuy0
toCNjU5l20O0ZxsTe1EHTDQPhMmLqIVuaQNcX8ENqo7LD6VIArK1kf5p6pzET3A+AEH4vDZWBg21
f+E+XcRdsenv7d7QwoXpB+iOBulNtUgAdqFdMO7anH46YS3KKkinAMaA71F/7fPCxKOCQngK6Mq3
7ZEweR+AUOUn3Sqlv+aAvd7Dmy9y0E1jMW4nBpg5sTroO8eK0XlkZyU4Btzooc0l0zOOGPQ0VKfJ
LOP8hMrEkpfcnz2LHARPu3LayIEhLNqd3V+m5qXQglX4jdROXjsgqDPcdS2Dmic7tqSkas4eAQbF
jxufpCdReuKmYkgG9OXZ5IIuG//EheFBUTzzvQlcjkgXuipuZT0dwi57K3QXEoLatTgp/MCgsZwp
RUUdC90bTS7bNoxg51jf/LvzCXtU3+v4uM/vAQOHrgJCYkp7wzzQ+8twKQK4ds4FXy+1LiW+W6ng
/EWjZ2MOGNgAxbykBwmGuM1g6tCIiPM2nb2YX8aikhjSYp4p90pA0ubbszigwEny2DYJxYg4qAY9
zvPfu2law5e3AYPxVFu0OdDbARCrKs6H/46q8bbIdtB8TKZMQ2dEdMgqTU7KfUKNSLnkCNpIROi5
WoShjmXMIluRFFbpn9tRS3umqelXq2NkHnre4nU3l8groO/gdmSyRAXQEO0U2uq4/UV1igCInKwr
/v2FOmPjTICIEKbvWkzg30qgvnP2rHyU+AbvVAzLT+hiGHbLt7G39GlAe0918Sa0tvJiKoORHWJC
HBzVsVkDg6dDATDtnk7JdStbIla4QsTsU4fo1mEtNb8xqQFZSwgHNVcQ23dBtUxihw3YZG1N2n5k
lOXebVQd7If0ky9xz1CBLhzPYmwYniqEUlGmOhRByBvQJ7FWA9nhwdgOuVtcxSS1/8/oLIvoQshd
EpO4mHmCKPapZuK41sdyvXqV/aUfnMMSOV13JYaVfSlqpjw9BQg/CMFWRCIAlASU1jCDVmIW8zxd
8P26oG3fbjhd24ywIMAiwrE0xfu+G+QCcDDJTWMzURO9oWOLEhUJUq44NlDyfrqzxpI+TYsQIH1v
D3/25tHLfnDEX2BmZmNG72NSOLu2+JN/Ozq9ECpd6U0c7hjmIFJZ6X0th4oe7A+kZToVcTmMykSx
DCaU088qs+F9IyUq5AgUCFJx1ywR4C2W7XwCWiIEWeenFsSi4fssP3DEURHnvQBgcRToObi49nu3
ZrgwVYFj/kpy3q8JqwF4mD0oTAZJtNRQ+zWyX12jQMaaHfhrZvh4sW9iX5T5ZPwi9QyoD6Fgb/md
dBBrJ6FFt/9r9VbH/J2WVYnaK7bYI6BR7HQ4dj4GoUCKtEj8cS6PLG1ZCUua9pE7R6se7fFfVBog
ZQ1RZrz4XV0ySa9+CuqNt3jVSrrlsY4/pqWDZpoksqoUsV0BXfQYpwKG50TiqW39Bx53w7FkQYK/
/aUSe6EVe94xhi1G/O3nOvoZ3+2hBqcW020tFwHNtFlg2U/rfCYqEUtyKUWD5aTgrEEembNdQcoA
6mDWzAcfJWfd6rkaacMkEgFLWbOTgufbcqoQQUoeJXtTK7DZKgxuI16Mc5Tolt1SrpDTJHv/fpxZ
5+F/UNFbRbRUXbCsbuOx6Ihq8YMLSyNKmNbRsXtyfVFwdEluOtc8YQSRI24CwWexpfEo1xcIMLFY
QLYPqDA1p5b+PVzfky4hzCor+3YTFe6gLFOop2x3GuFKyk9UXqv1OpYRmqXDUWRzyScfxnOFL7Xp
JL2stkuiIvPI7GXjLo1Y2+uneZgdPhdtwRLBernxJjCO9xs57WNKGfiyEubz1HRpBDHYecV5inXN
4lEzLAXYzuBQxHP3hizXAhxXH2s2HwBusaXXqo+us2u5X+jXZNneoLf6IshXaIchBsGtLyQ/JQMG
rn3WSPmOTADztsWnszLChborRCPL5EmSqGTuu6Sm0jJ1ZohU19AB7dbe22gh3U+etVmj6Fz7gBVh
jvyViUeNFBj9XA96mv3KpNB02GFoVIp3orD+p/ppZAPzUdFhFtTCuRnwgmPfJ6/2YZNQnetvJ+VR
Xq/ewKyGOm0NSRuGNeoA6K6ex9yINc3mXv5VwOesPViqGDwIaGl9EShvB1ub3SQKxYuOsE+b0Gct
I8d5CpE/O5V+2ipoAOT4TMNsyn7RWPbZSyk1QY5Ic0tL+Mdd3RdGqcbGJxZiwpZNoVnFypUywyw2
301IxM574dwIfuBGM4XhrDvCMH8/cI8D8exrsHaF2NRb5YF1D4Qaz3qJpEwbb/+9uEat5PCQBUM4
qOxnDuk18Q9gz3g6X5isVs78xlLJBvdYJAMr+Z268EWhJ17F5e8rn6lzRUn6z8SagFBFDQjQdT/C
wt7GgV0fNJyKiiThFhhbUiQbXmk/+8l7NRlq/et/Ah5eIkiDyXei/6uzvhXIActHgxU4IUl3d8aZ
irMh/8VNPmaidGXwTI9EoJKXxjansRvehBR3YExfKcIh8OKd4lWZc3PfR5SjYdknwi44p6auYOj4
vAin/zal1BF3BuLSEE6j2+42225KwVRA3IjUSL+BrWKeI8Rl9jeGfJII2kbao2Uqfsi03lDKPk+g
VeUDJF9HCPry67zVvWmBKA4pITQuZ/PNCT90T1EGLeDFuDSuBievl/aMJKhR7UdOCJcmGv8vSFHJ
zNaSpqa1ePYg3GBeRRbXTQe07OA1P22cv7BYPr7CJnQHogRK+lbAup5hr0iLGyL2mKV2QkGGv8RK
CvHXgZEMYnEIrZNnund6YZj7Jmr5A8DdOiRNbUqS7UW5fFvvmbo/yBTPyxKwOZYbr7Jd8B/h/5O1
dRaBkhnGhNfa5DZ0y0OWFSZBa1Kwc4jtqxB+Ahn5EpV1dUovGinXc8CSdjhwumjt8BaWRtdsJWtZ
oIuL2iHFU1j1cCqGMQ2Rb2By+B4rm3bREw4e5aApWaRtUya8Z+S/TocCbA6lDyA6mQ7Ww4NxvVHs
enjuducLeIOUpP5x4FrpoexhjdlLxLGhsXDaF8bz6jrqPXbByMWSmByBU9ViZVH9TbkSdWBZh97q
Igp5/rDG0ak/23XrUU5iCkgX+nk0zCs3eNOzSrT64v6Cj/MHnJzxh/VYv1bWbmrctE1VYSoAKn4M
xgWfK7gM3y1RkusOFtkyJoIkJTIrmK2mxGyGB/nA4ucgM3J2KZjdCKmVrNkX7QFZlf+uTUYwQqUE
pneNPmPK0U5BA8H64yBM+lJ7bFKvNeSn9ohzRLMU/HzYPa4oqQUfAiW+WaVnh2r9PIG0IX7laiD5
en+pAl0eMN/SYTjRw0mEQ6yLcfLGPc7VlmOKQRAP4mJkZtlxlB5/drRhbEkZT2MqOdqENz/42Xzx
itaDpCAI3eNbevFcJuhl7kVlEB+yBlcWfjTjjLOVtKC6Tj68c5peb3H2LEUd8ek5T9I7hnkTUiGK
B79wE/2wLtNINm9kMgklaLg/oBfNupfGXe1mbb499K2DsYkNBKwqGSTxuafWfWtebbyqqZqedal4
EmbpxrVCWwGnRA2ntJL93P6Vf6iZzpAGo6/LjSoNIFIOnVbdn/o7Lal2jC3Itg49B1EXWbAD2RBi
QMbb0tO/PRHOrt4XoyfznqgO0KxDC1y+Axa9/DYpUxRFqS9pin/hIW6Xacg9cSWWmKih/szwXeS5
ZNx81HoynnqLmP2q4OLsj8k5q2++AhnFP6ovSHOFV/ScrWiGDYm3cuJPLU4uazfdn6A72gQXXgMZ
3q3ioteVuVZRIsTx4ZLt0aRtfWygh0fKWBr3Dld01FYtthZwEDJTCoQLbBvprw8Q2X66Ja4cXf3v
mLmhTutAfxwHQH8MMxm+VRGn7CWsoB5D6JaUC8DrONEgNZ3tUFD1fm0OLmmNfTFCvZG5LHLsHFLf
OPUPG9pr1u3f5ybBWHCDkdT2FjW/fw01/Kc1Auilh9nr1rB/7UUO30AusVtQE5xJenA0vF9QtlqN
RBNl1srEcYFpF/BS1HQbLfbqOtpNcPOlGHPoUfO72mrrOjz5bOYBl9L2CSFze9D7e2+xnNgIw05R
vHe2fTPnkkeA2Cz3tZ+Kd+UEOs36qjW+ycgh6CSebhgw5tunD046uMeuujwgh7eQLcVynqyjAg6q
JQ84hxbfW+WiiXYPfbM6hYKpE140ZEWUZgmCe3ivTF776OGmND00MZnZNaFoEA1mjwIeqtub6ToO
ac1ve5iRRTtnAnFAZzBoxzEtt+CozDG4ed58sBbmpQXt+6q+0d03Dw0lHtwLJkRThlWsXTxooEt+
N1ak8ZUMcKIH8+bQut+IW8h1IZHF01c+LrduPMnbF5Vwk3xpt2W8HNw2K1+v9B2QZUdVduDy3ZRq
ivOPnwk43k5P7zc8rVSyT8CTymNmCbdjFezjqJUFrbdVvl6v8uxou1H1wiXklYtWS5yFrt1OxzRE
jPfEuXQh2FEZ8UFtpy74aTb5FU12KgC9aJ/p+BMp4BJI03rx+gUNraqq+tBYFXU08rW1iQZHVvL2
Tl+TurIyVMYaAcH/465N5JOkLJsssrMNaWMbPBGtdwULjiOQlycURB1KkCNShzMH2s/BiUcztDHV
3U2/RJ6vhJRzlQXGRjneBvddtb0cBLMfIKkoJZ1UvZDy68NCc996iFYtSBZFjczi+UUlxsNQ++j+
0wBcaPx3mdbbE0yQVrF/vCPbA6v5l9h/gSzmN3DXK2cFGJo1lR5/ZLxG1rtaTdY0LuneD0KweHRz
wcu5R/rAEsn/XPxY8e94x6u+fCrQpQn1FcEsWloJ6tDiXY4hYy3R7QecAFUZfFjJK9PDupjgbHwz
Nx24Oaf/7kwx9Wx//PFd94/QXpqXtuKQfQ0QWTVBvOKVEppRQ95CNdhvN00g6XFoVFbRWp8X7ssB
Y8vJzPokMNbMNbXm4JfF5uc5EaN6afVHP/d4zn3sCEftRnwd4pQqqdqZz1OFzYuh1+q28nYhlN6p
w03oIZ5GjReeA29562UtarwImQxScWUNfySHcr9lQqpjhIudpvs8yLfRwT1cNp7mRxgSA/zeHrkM
fw6B+p8YLQCnvxuvQUnOH8bohw6MauGReuWDZ/ngzNGAP7Im363ueaGHpT12fCvvwmSVq4Hxq7cY
hzQVJR/DHlEjKbKjGSKyoMyX10N8I1tUfW3XrakJq916i/uVOl95khvA6bbS1DwaSJHaA1BK08KO
VSAHlZnSdkqfYnGQyaM7DpBrO63wH2MdBOVisKDNSg1inIXMPk6keb7Vhfhl3KVujymWsS6vZixb
0Fnlctm89KJspWjnteIlDafxjqxMxOo8sL39wYqOiSxI+s/J+ms0qQLxrdUjLx7HvXhxInEO/Dpc
N/UpfgAzqfFK461Ha8YL37KiQPN+dtRZNSEEB/a+mm9ZDkUje8kv3UAHYfr9eVcU33UrunRHynaT
ZWiUTkAFQVzaTk05Z4Bie8NX3rRJE9gjFdIVdh/5wNuN71Kp/axMu5KUbPPSlpzA6h7IgtG7sMMp
klyOCcY3Q47Q0cuoFFN+OodIxU3RyiQHynPfSzNdzwKL+TNAUM1Bmue2CFqimYzKb0czo7sB7G35
tR6y3DzaTItNNODEZLhkUtuiPSHx89bmwvuJ6WiDAfKZFMlB3dmMcO8WNI3h9+d2W04GcVvovbKs
oc8XmEO7FyD+xbFjh+MZFRMJlTQ6s9mNLXoAdtuC8CcnmK/f04vVt5BkdDusW2hX/OO48a1KyAsW
erM6/f2gYc5xtpo/I9eMG5RmUBvYnO2+vX88hj+rv04FepQdEJ1XUE4ClsPrt/FuZ0l23IQgLLbh
5RGHGVSTcNGrAuowXJl9ytHq083TDJ7dmGqYsW3ZOvRF5SR5frMeqXvxuwCdLq0cDzM/Ta/XJEjb
TKw0xaXAS1z2c1kmAUgqYcL52All2tmklWvkPo8f2A9Dv7qKALtpL15R/XwhjYf8T2WhuWqSVFW9
p/yb/oZxZ9VNGHXD/ib0KOZ0mcymlTw0iLCh8lEiMhLJcEBig3GPf6lXspViiWvdDne8vQeX12u/
49iXDlDTmQVsNTMrICpZJM2RcjHjlrlpHvfMN8AomK6jA2Y0QxnNv8IT3qhYsRFPEpuLlJr/9Fxr
FsVLzYp52F/tlJyuZudokbXOltm8gq/tu6kDbTLgrm071IH9wOdtYgDV9tS5J9sN9Df2wJ9E5Nzx
t8GiP+zuz1YTa6WXkx6URQWv4R+2Ov9OJLT0542TcTdI+DrgL+sIVu9feY+T4n7qhiER60ANhlgg
cltSj63rtUonXR+dzpWymwzZkMZsYijoC1xqhker9PPhpezckKJp2dY6GBCpc+rzOxUaDz90sANn
ndzL2/1y0ROffKakb/nZwrkq5/6eFuxEqXIjA5obQSknyGeNmRIvS4zm9sWyd6xghd/aJIZc3OlD
hihG45xjsvnkVOTckJEZDRQB7x4YK/VBCaFKURY9TVwuYWe2aPQNOGRJK58YB3xoJ6rZQGgmI65s
E0+GAjfmrhqPTBniLxQ1sNs0fS5NvcFwxfAyUotGNjJfvBr0OWoj4sjjP80Zg8LigZOQ/IQETN9/
UjSe+TDPYPQbHZPer24gCkfAmGeX9gXhYKrE92oQ60L9WXsW+gm7I10yDv6EdfSpbxE5qgHDpz0S
QLt3YmzBCi8ifhlpvsh8APwbDvD3mtHq7ydb58pwKYytzhlz8LTz3Hr0GiKFWzlhSRuTDXHfPVZb
sE7HNZnmmU/JVBXLJEW39nraiZxTEnEu1322RblKPci1+8FrFuPnJpogI79/jPYSSmmfR3SGZfml
bTLCX0BDRGXfdwzxPZigPfvYTEDOkEXRo40wOojlx+sr1HvUuuOer714crCvDwJeXiMtBGPB8Oqk
bqVbJtCaPDaFZ4EKr6ajGL/eaxe/1UOaKE1LHUMoLS5cUu0Ozm2/5MidLTy2nsV6RZ7pV1a9tSot
C+DUTCwzRK/uIY+SaffdWe6i+ZIR7GHDrNmzLpdextvykPm6u9FMSZGsnHORC1GaUWYVtgHdyUl1
dOvIxvnuQTHRazdrMAxaqOwl7E2cCzFN5UsbfH4sSO5UCOV3hF9lHKWB0vwsmEnSonIuNDet/2dN
x4bsetv2K/IySHB6qVIBC/by1hctq+qmMRNatEf5HzsGzOpjVrQVwQaOrqoqu58xdBHTNcqp57q+
ymbScVt/pV2lUNmSEggAKbzXEVpsNUb3esKylIXw7SA07sPf13QnzIPxlOR6CvGUE05uN671YHwr
pkhDbayXyvrBEHHmm7x/hVSCs/2wJ8pa9wYlvTdnmEb9Ae+TrAYDh9rBsuUr6PDmaVclprkdODI2
MG62GSzo+4tkFHYIagxYn9vE36G/RS78AQvYbvdXrxFdcLAdMqK4VffsLC2NH/lgKJ22SskKuk1x
Ek6b+m4fSa7HXYB8Ar1SavPTEUi7QdHxWnuil28RYr+2UR06KqTlOSJjnJi3n2kYRTbigzA179Pw
r4tE6oJuDNj2XPzdqM4dlcvSR1Ib04HEx6gAYXO4zZqC+dbbEZq6DbKeg3IGZ/EJqY8Q9UK9an9i
jLdG7rmU2Td+zfzTlyD272AtAayxxRjXF6PRgb75JIv2bF60mJ+VXip2dzfeWwjXEJtVV184bkJD
iOKu5OB3+PsXgolFTm3JYvW27WJMITnRckgpOXi64BwmgtVCap/df+dg7rcS/gDAiAy5vVreUp51
3RJj+PGMBBcLap4MWw7WRG6Nw2pwp1Kr5l1dO1lc6pkyYEWReYbiSc+5+w1GmCl2uQWLJ24hhUkw
uQpJbGsKxpEHITDfuXp1UUaz0vsEjLPMaZCja5fBq+6IcIQHkBFYMp7g1ou59JajEVBO8bJBLdsV
cB1a2iqG1pEhM6XJ10H+x5fI5Ym1sK5qn2gUdiJxcC6J02K0MGfvpJvl4X0ZmqeG5KsPS7YF/Vt2
9xt1vdKwS1Y7095OL78NmDgeGZZvcbHSEMRx1VoG8es+HtM1dYfInYnIUHe6iE/iQLomcO0dDzDG
aoAj+/32Zauw8K+mRq3qT5BmzPhD/GfXZsynclue0Q/QZ0SJQqwbtbdgHKKbIIAMMQ9V9P5O/X7s
7HbCDNsaMy0nd/lGQ0f4Eafch7b78BgSK3kmtD3l8WYlQ9p7f9dw/BnfCcfe5xIa4E19WQDOY+kj
K24foN2py8R2lresGYx3EG+3UpsfrCD7f8ZdJNY0cCbh632NsZt5JoIQ+st5jNyW4A8eeqUekDll
Xy7TAgi21cZDcgk9yVIL+v4KXVGX2OXYLbP02/bOR8444VjYGxiTdzY+YpQtZ9sU7EBs+ZW2V0kT
v85/BuUexwlhSppGzkrjiP+jEA/70mdffG1+a7q4K0fZVZ0y0GfWzB4XqB4gtnvR15aHTQMl26Fx
rhmAnsMzVIYB73pDXCxP47BcJWiMegIk+sFozUbWm+7nYj92TUb+xzr+qEaBma85/TD9jiWQIfPq
Hzhd3FKc75/gDfTnC7pFPp62wHTdOUnf+Jhgl4/ELFBVs1aJ2kXoLBu/E9GdF9TAoM9eDMb/256R
Hx05kd9uUE3YflN1Atg4Y6JEFfA+O2I9f2CPV+ZMmRyb0CA8YUTN1ybK79PO5ey93yhgF7Q5AhYN
9KivoRq25pFmtuZDBwA9WXKyWjVAQhcyGtYvAt20BPMLn460sW40h+E0wiT/qLLO5YApLirDLWFz
26px6QpAUMQCEG9/7O4WWKpnIJgBIvDE+dBZNfFvvCtkGpJrKhJif28esbIwN+xtvxGGvLqSmD1q
M8pnBmEbd2tyIGVnwDm41ixXGc7fvYAttNfYoftX8sR4in0SJ4iA9LQ16a72XZbkbCRzXxJzmEW0
5YVrRBlB1YflxqHAgc7wSLh7YV03sN9hgsl6OwQexgnyShZXBbkYaPJfQiQbvjSPlV0mVD6a0i8G
xAIjV1yKv+fa4mRxI8B+B9zWHzCm0cEtuPU8mOSSA87n16LYSOcGYz6x+T3iROHu/bElpeZ7sYU9
VXGpBWNtOjQVlNdUOGUUUDxs4G8ZJ4bXXXlfd3ImeyyOtVxt+eZ5hVEFXUnS18APs/Sp+7zVE7IR
fIIHR+3K5qnB+1E70SSAEbwOK+1yRNYIaCzWN1VtiOofAHvwiCQ/aNDvA5rHJVcwzfqLiA/6nsTz
cV9zrXpC7bO45ANq/2Ab4eKd89IcSWsicR2CJHSTv00zhUNTUv+czSG1xJrLuRihK7XS5fOo5u23
omhvz4lkjROjz8K+JuOuJxIKtZSrikvzh33rrsvfAxC0hBxPXIs9l1ENNtv/VyfoNsFjarZrTK2a
4Sr5n4NFP+brCx8qBEIsEyJXxmApZE1mP7YN58BbR+Urh4Gbm8l6F9cKyfBQOj5v80iWnOEPsnS2
XgmPmmuQed4alOhqTI46+MM/VHYP4NjegBl3Q4FPIqeeE0LDFe21AOMcW0PmMFHl9d2csDD+RJBS
lI7qbRQgRkerNGFVf8/bt3hBLkICzcSkfH/6WcUhDlnWiIiBS4HUXSXnHbWvySBrAy9JvsEKeIV7
ZCSTvLK1T173Y6yuvH+mpWrfeWVUYA4HRqduIFcR8/XGSyzJG1CxcN7oFIjRbj1IkKz+VUB53sEQ
NhQJpiTr2VM7cjHmU2LNNGRN7cgplpSCNEiT8ZlpRy5Sk/UzOdqWbdEUQXVuTx+yB3i73ZJrfH1Z
hERKeZgDR0zjGyxfwJc06TP1JijpozgPVIrgSz6Ga2bUpN4Jmnw32HWGiQpgT5i8Htl9GKaZpQmA
KIFOhunyliWcCf2RKuqmvLisTcYkvS//EW4+0N233kakcrrFQA4DnciXJEOk4qGn0UJark2yJ2jp
p6gFOPqDZR2rwHXtwJZeSpfeaaLnSYy+wDhvWEqglpdbDUeyQxw1UkZAlrIbpBxH1XL9B2KT2DhS
yOzh0gvFoES1X/aTAJb4O/6hdegeXg0HkWL/OZk3LZHueYFATud3qBCwYeKnZoKWVozs2EvkTsii
ToY2cINKg+dg4cn+6O4WchXlPy1ZAmOcrVKtsc2fKVNtjVWDaCPvB8m1eDW7CBgqc+Oone/mUbip
+jsejW0rXiiiQfavwzoOymxG5uJHDKUuQ1VVYT/k/AEpV12HGls9oSx8svjAPzyB81FXYgJt2H/e
bKzPtZGcljCFoIKqhtLSD94rW9QM8JmjQDpIjhq1C3gW+ilbB+0rbZqJP9+Asb2mtiMhjKajjOC9
O5+LrZpEL18ek7+NiLC/mTiRd2igkRj+0UAbJeyjxC8H8yzTW5zXcBLofjJpwL0o6X9eDsenD9hw
U9jnOeYrMl0hU6LyI5NZ99LkqEC496bEphbjQexJtUkG/7g1Sv2F8wGRgLGUVM2cbe2dhhi0hck6
9o1+XWKnh5cd4jiYHUTP9f6g0ZOLBdKAKn7B5i5yl535Hd9otYmBwB9Kxz0IXvl/scNn/DlXgOq1
ivoo1rDFzM7TGcOzsgmQK+3Hm/ddVI8Ndkqmz9353yltQ8wnoZPC2bV+zuaIjF2I4R0ASZLzQzXX
LZMZmdKC8egi3czyBpergA8bXr7VjWLdt6zxrxwjbxHr618T2CBBDPsA/e+bc2ZrdgkRYARaRsPZ
+WzY1quelajSRze897z1oeBW0H1e3zXLQwFapiFcU6stDnWpUd53g5nFiDIwSleXN8doE0wveOyr
8S5TWcx/3qzoin+4MqKEGdQLr0kr29YGGV578v7QNf8f1trCJgQol18cWSKHXb25UFEz1UmFnBKz
xUbAIzAFDWnpytwLkqlehkKUjAU8FhgwvsYimX6jQ9P/lIE8GA894BC7AbfvTKTQvTxYm3xrsmhL
tTggIAvK5xUlE5ZMofIfQGYSeWsTeKHiCT6tPCO5oYJhPKOeXnn9U7H6JMa1M3FHjJkfqpRub10o
fo3tr3YGFUmMmNEwJKmDq9JqL/qRd8XbWDZDiI67oT0RCljpGRK9JWkVSSvg0e7ZEFGKyKa6nnHR
XSMttdvV9+nM/6BVE7gLNR8nlTqfxzBOr9jqEjQbaMomdtIqpfRCRfooPyQAgvaVAK0JBzqIDf+B
7Y5l8H4dRGnSZfaIQu82Oo54qrRqiXMjvCZcXbQMEfDFiNwMIogiYleaJv6o09DIck9sBu3UibPc
wObuw753JCtlqGeRz/pZldWq7scW4mZ8PwRTYEImHPg2mFZGnNpe/5JbntxA2mNbrA1DKnwbBqBk
+M7JITy3OcBAGNyPNuLhS7qGZLlHdZ2Zgpkcj3lSGLeUsQ0sjkATflkdKN2sbL1EjHxxAoX1UvFW
adQPjA4Wia/JHYR6NJR4sf2Tsvo2y1SNtxVYE0aiA1o0z9/hYO/dLPUlVeLWxEHh/UDzQ7UrYONX
oBudplrG9rQyIQrAJxUpq12FkYi7/0f6GVHkTdotcOebh+jYGsIy03wLbXtvpjeLmzJturrLKHBw
5e3hvJGyPgox1alvL6o/ZE7Fn8ADFtuog3RrGjuy1e9eE1r0sTFIS2IO/6jga1jnzLK5TQp1340h
nWd3xsaXBRzczSIa980aUn1sUkBcMUHxqyZQ8Khsamfid5I8pp/BWlNjbaDlTAdo7SsBb+2rTKPb
kdwFHB08qFVA5CsSkYR9q1CEDHWDNMC/P+HmdAMrQyQAEIWrM0LUZAsIs/MSxPk1GhsiUJwRdWmK
eGhNXEBKXRMKzlGmNKCcu8wMdy4cYnabxGDzX6/Y0buTwuHLNqAWTsxe4YrLcCAV9+ht5nyKctx5
wrn9tGlnUkM5sYDzPDS/7kfzUu0eXodNgwNn3sC4i7XIh031BCRW5Tz6/Fu5GNpthijQmrIDlDl7
RRDOGD8jYRbIbcSaICRQVyWdNo3TGpg2ztdXYRMiBlBN/Vgv3V7yXHcDjy3CSxP+Kz/jsMw9KYU4
olXXlX+hdRdD8+/A5A032SKNyij/nI9nawrzaog8+20HzRy7+5aMSpG1DvjfqY6SOuiYBzrfh9+i
Cn2nAhiOQoLw98XgNFP3VHwWWDxzWJIPMLwKpzKLBHz2zsgy7r3krzuIY+Y+Va9rMUPoN5D9yNtF
/5GN+kWh1aSGHgc3VzF/l1JPueYQQRDa59PtWKU0WG0XbCo1dSYTgLWK30l/KnUy5eic1Bw4cvEe
chPXgriAJNlyzDQf4tN7XElNQ38GhIV96WnX4E5gsfKEkzP+mKNXTn6c5VTCs6p1u3ih03grx0SU
JCNVuzNFF4MMxUL3qGGUvIgQUraPjdTmOFQvS2Nl+Xtf+IcGW/aTkfNy2UM1/VJrwCamUBYepc+7
+OMczRP+wh4nC1pUKPwUKpDOrpCXCAPWJo6dKKcvNPPNat05l00i2Mn2hOsVucJZrUkhTwkbjbpH
b+6Oe2wExrp/i/z6a66+H7z29KCU7xlQcjOty1hcNZuBzj1e4yNXJiiS/WNW82K4xMa+ioqHP+0x
LBKBu68O+Cl44kv+ZooU5aPmEIdJFWQ5F5DeC+fn/4sWGD6bn9miVIaswk4DKe5QioJ6vJBDRXio
/MrJ8SJNTonzzdTCGFAPbUcvRUsf/rnsunyWnad6ysJdmhKVrm1OZaOh89CfjVEJFylZMvD61m9J
deSIEh+3vVFNGnTgbejAJF9u71MYmCIERQTeLzLVFO7V+GcDnPhRyvQEINIFKl+iEzBu4DNQD9Wm
gG7XcNbYioHZ+A+ZaOilLs1uSGx5Lt9f9ldZraTVodLbpvc1pH1HZnnkUmMu7/KFgBKYFDYmmd2k
DkW2XIhahCeDnrl0r8KdgwQkq1fE+wSW5Z+1BSKRrH889lqnc8rBsCrFII7HxkJvULLVwfSRIBPc
9aIOtzg848KUnXFAOuVKkmyGghyqbIhDcZAondmDy6dMM1blcICiFYt0UqIxVFLEFiFFwxyui+fY
TWeoOCzAa4CKu6gl1+a4kuAvYm5coQtwG6hIgaz7ROnFZ8gnfhBFW7CAcPH5kNB1BLYrzf/AAKi7
BI7JG0Ux1lgCOtGCnPyMGTSI3EkktLUm4TeLR/+jRn/R+zhtP3niCGopK/RRk4d/RdU2/oZa7wfR
+C0If/1mmE1ri1Y+cKD5mE+I+vgFsiKvvg1x6lqn5PpRZp1aFakwK4IaaPM1EI9V1TsLk/y+FG3i
TutWXUmQtlStf43CLP/grpL1pJjGr2C+hZxR/RDYJos3+izPHhSsbdpU6rArLdcicKJ4YlAZGkYe
6kh9KPrBbNphi+9uQXglHM7q79Hx6/CJdUdyOMxGc9fqp8bI5K6i7RQzi8X38aHa51/UI3Kuwqoi
4aBDFx1NGkLpq7oEjV+754b/MD38Bgan21JkJZ+Yd107iNuZOM7pYr7cizOvLKlNOHofI6i7lUgN
5A43r2RXYU/qE9Yjm5HleITsVxvoBmnxtAAqWlRDcJpmRRf/6jseeflneeQ6ZsRafzcfXN+iPdiM
DcUeeD8EXuI0JmOMbMw2SHyG4m3/QUEMnUwOcBhe0zLDNpoxOMgyQ+YIy2D37eQzd/sLQIQQT9tu
pwLeMyOqvcaKLrYzRBkzOjwNMByRStvM/wj0+Kvhj27NckK0bSmqDAROB66cDFbaq4M5bzPnohOM
h0Pf57PghtljAcgsPD4YIMWbhMvCBk4xrqhQhLyASrVBpPUzO1nxWb+iwMgDgsSdO7DlpluGmE5t
2o3CSDbrSIYW4jhKJT8EA6/epUpbQMk4ESD0KBKm+tRoAUCF3V9Nu6GNXU0yQwg9QDOPMy/FRa+o
twz16b66Y/euqUD4gEcXNsA1CUeMm7YzCENIfWHwiFFO4dlZEMby/p96zPz4V4k9/ojGKy9CVB8x
5cEsSKeuKjDXHyPNSyp2+T2YkW06jxGbAF1TrJKge5zS18VZDwBFFQ9rcJnB5PfoIvMO75SHagT8
s+3CfDv4lWTkN05WL81iAO/70OSjpGA8iC/2YcQKkZZjlF8MlKYrIvHiNACNcvtrL8EH1A56kaaX
4dFwFFJYmOjGXyllOS0vt/NWvImQXjUZUmR3S0Xbof6A4Tv6SYYWhJd94qJglgWE9fcvF8d+Sdqq
DogZq9ml1QH02zwFYQeIdHFacQWgdvDX7xb/oeilhvIlZ+5X+FRu4jYsgy7V0X+tTGflvZKaD3Vj
GtatSlt4is7P4lgvexNQ8V8Oefk3V+P1YWBbeqVGSpi9ZURk5QHGqVG7wR6sN3R5W2G4C2D+ikp3
G049c7tL1hwzjPNUs+YNT6FZnPeSTlnIMsS/kk7VALDj3E9GrHTQyq9zitG7uuKjVWQn1ShCF+WB
oPloIFKBfxRDZCHpIZx50guBes3BzlhN9naMD28mVT6FhvgY+abDtXnCRe1uO2O5TEr/uOmIRvRF
9XsoPI/zgP15hLCTIscWr704URBduOOEtJuaQM1OK2UF/DcW9pp290dE3i9+kr3G/1N6J9EsWxWo
nT14kn4v5TblsA0InuerCtfR91JSNWJGV3cJLn3jsP/U4wB+7lFlvK8h7BD87thurcoR6z6k5f3v
Pnpz2A4+Nq20MzcFkXFf66gSChUT89O7ynpxFCsiQnwr5JiYdJH4I6W2GqQCdoi87UlgG2CHdS9M
T9AWaf4hlvXbrKR+lK7BOWQ/CzyDxtVgXIyGsaX4S1iWkt2GjK2nADofdmcQMF+qjMQEGtnIUf3q
wal8n0insfC3Bhdnje0kKrTAdy60caka7WwlUMRvl2q0jh2eTljK+b6hoysbUd/6RoST9ivgB4KH
cDT2EFjUmZYyI8aC7tr/zltTup92vA+zI0GhnYR83xFoHhMXkLmO+FeI/zt4S7VSyz4VKKMZ0BCz
vbo7hJe/DjqFdUPl79V/t4MyVLw4/m5WKwf/Pvp3OJH2RPay6/AcJyJtm/4sKsfN8U+REAXmCJRi
0/i9PT9bTtWu8jkuAXI4ZgUF+biiRZD+GAngEXZOjUGPCD3MitbZpN77a/VMwtgwkNBmiciHHttc
uJhENiP1oeW+vwb/6+yEviTa+0eCFLUJQsvKmz6uOnR7kQvaLnfv3yG04Dyoc0DUysLArdAQAIBN
O3kmflaClXxIr/wrPPHkng8bG+qH03H8lBURfRuS4hRoMGNto4/4bVVkq54Ja9emowWjNcHqjIxE
mfN7iioucOg+YXUR1EC6VcDxDIk0Txlkww4WHGIb/5aih9f5KqVDtHjLqCAJaetUjA5YH6PjmCjh
oRHloSg+2AYeL7NEupKoj9QZV5PKNRx7ruxnLdl6mT03WK/qevnaf/+6S9YhyiDh60nQPDxIkMh4
lkq5WA5KwUll/vvV7z6vhOP6NqNKw47Z5fpfPlQJ3qpNVAcgyPScALroig2UaJ3XgQlxUcO5y1WR
QqcH/qhZ//qqngWNgZriKWyFTZfbKzquRLvFJMPNs5dUV5zY8k85GQSD+cSkWodSO7XDf3+Fczy1
8G88x5mXLS8f64MMg7d6JFC57tudnSSIl7jM4X6lgiLKDLGoyNFdEYJpKBhraX9+qF+ZYcHcBX05
hAHjqEeqJMOy9GqDS/0ggWw6S0s5On7isKiA7XXwU6Nks1PyHemx1Q/JpPm/byVdCRl+92YqwY+V
5H/j4RaAad3s+mnRil6Y14kN4BmUAxndKoXAeGz2v1ok8DrUBzIKwueeZyVFe02waqtxUYafEnXk
TKICKTVGSkxfnCsddTObu26rK0QUeFvmzB8tNyNVUG4HB3jk69MdR9OuqB4Om3RmuegzksMYzxdq
RuDPFEHilSmxU1dWNJwJYicA4sSb8tPQRUAM2i4OMmGiYpX7PV8tba36BB7jBxDYVp19/4vYUss9
EQy8TBmXHE1rb24CqFrkaUrCDhGRIgeImxLXT4T4SIt6tBLUUDKz00wEN3r8knLCEipQVPIBj4xO
kUGeDY4iuA85KPzcHtTd3L4GEU7e5H7RAdsVK19q2qLRefVBv0LBfLojVRuDRvTfdqCxT0wL9Qxw
C1MDTzu4kfoh6saw5RJF90SfUbTtgl/xttgNkciQ7+yfiD9U5IVeLZR5gr94bYyIRXMW2KnCDCfv
RrKOYDoXZN2Rp/TQf7EhDoh1MUybtJW4j5TLURQ7rwNtvcT5Tf+dlywy0BfdGncf9awJtt2b8iwc
n8exVg6iIRAB3tD82SRh7zzaAeEbzrj8jdPTvcj8qlOfXNAtEJy4IXP9b0FVPW//7b2K/zqLnR4W
w9b7K0d2mircbNhjLAqKqZbJZtQTlougDYMZMyxlcYULIP1NCnKsuBQn2m2BQ8aBq8WcoSrNi2lW
KZlyHUlfMOgCuTKBcM4aDdq4yHCGtgrzexO2Vw+IqnfDNpl0FrrkQA0Nm7Pvk9cJ9Zqb7kUDRkNP
35xJeoHvUOA0sPO9znGMn2zgJDR+nqcoWyyI5zNmaBluTbQM/NpQRvkK+aF8SI0muqEy7KHMZUxf
OC0qmNdNsYAiih6uqzFRYy1BKrfEQpaznqhY0mUg3uzhfEB8I2Xll/0yoVLl2UZIliOKo0jN3UnU
qD7/o8ED3pHsRq6rhod1/qSuARFpTFpkvQtIc5ZywLsNHNsRp5dUMSc4IaA12HW58ZZOi4T532wR
pndGAou8wan7OguxAuN6sDbdsFK4KElnJ6z+Dk2GVOQEi1gP2Qky2t+vJxkzz0oAom7jCUoBo0Ik
3ey/d2TxOpd15wsj3B8Lo78MSVXdYMCsVP7Qm7KwWCbehFRyT74CaegkSPvGmgI2tMFL6J0myPB+
IBrZJF1MuSxk3xS6IxPkfqWbjAFBAlUnKC8olQPx1jZJyzW37KhzWFz1HKgV6CE4OLsd/gU9AQ+A
/uCn75s6fUMeo9j+THblr/PrGs81yI/DCX2Dx2L4EykdmoRuCi6q6cPkjmd1RJZ8r1mN9BaG6Pvu
uYVgoMC1pbAO2U5OxByxJjYRSRPSDtvUiuDpHzLt7GmGocvq/0PLFiV/il/cKH63cReE3Lnad4Y+
ZGSAY0kLi3ARuv6kG85kc6E1/qeg/pe5r70xDErc5slB+9R6/l8sAUg9EHnDhI8WXd6HCFThZXqa
vqSrV3Rb98YwBSfBvdGAt8KKqRl1r9igFrPPi5/2I4kyEgGi4rt4oHQs+HtdvG4KSGkWeG7AjoNw
WvTzAvcz2GhOOnnGESfjYHKisONAWf7DWYZG/GIrmxzomcPRK0REJTFr1HLo1X56imQKC11t9Bpa
0ylTIEbwssZd+X5SYss4p3cMloIt6CDBmQYPYfWj1uxyxr277AE1OjMjpWNLodzABpvwKDxTLPjf
VRCZ1QkUkJSome1VaRu/y3oOVZszW2KYmUzz9yEfFy00GldyxRGtnMznLdodfD9S0Zjds+m6dU/+
K1dDodmk1fqu5H9sldwMJXYcqgfNmrXhmL4B34MYQwRFRtINxfgVxKtH+fw6rVMAvVlaNH+psZ44
fypA4wYV4mm610Mc3/6Qpdh1i1tClH6KkI0zfR1HhtR2lrw5//VkjTmcoJlwq5qOaj8aJkC3/HvD
x/k5w08XJu+NRz2AAwutSOc+S42fn2czSoWfbEdvdNtFZum32iOmgiExn3sC2fyNI+7B8p4/geJJ
uNECK3126R7LQr7c3wvAsHeTT3Gi5niY3sESe2pQSkgSMwwFpvFLnxvCs930uvP5ZNQ7n1NF7zcT
tEaj/4X1M02KBroU2XnDaLrlJ6wTlPbsWWezksV17Uq1JfT+18P7Av6e3xaexaZ0dAUcTp6JTPvh
r3orf55wECxf6+5yVr5vwjMpyqzeDhLUclv1PSwrwngn1Ghd11bi4TRBHZl4zZZQbzZxtJizt2Xk
IE+f4NIQjI4Ry9y45lSMT0oGgArRUN/jCXVotZx40ByzooDXfbNbHxieGnaM75rMn7xjC9rEQg3+
e9+SNeDq5tRt5UdUbSI5JXcsUkcUKmbN/n8yhV9LB/t2ACoPl96KMEhfnD/kKyk/K675suoGVhMH
inNM3HD7ykvI4EZQsGmYgPjurFCRPVPO7Zo27sGGvtd8zHbtLZu4Lckd8NlQGDN7orhqytYwZq/Q
a1KS4KcKIJ9ccq2NSBNVH+lRjgbRmy0SYTKYV9SiplS59xdiFHA0ItVoOyfnsyEqsaw+TJ5W2XAC
RmKLFEMcAPYYBfY4gCJMglIwaTxjjq/v2+4/2Q/sHubUgQelVURj97uiZPt/DYVrJkntWko7yJL2
kHWQNW3A0ijwYxTOkZ8DJGSe4CtMAM1OZN5xYJoP1XAMJwoNQgVIyuo3dFQ19YuObvbls5ycLPAD
LGK/I0hCg0JqpxmP/6rJ/cvouD65OKhjJwqTvH1czy6X0MN1y1pJlLKnvEzhRu3peJ2yCCe1HZEr
/Yvugg63A9blGkPuwDqIjxNIIJgty0dLf1t5XgVgPeQdMJ9ZoFV6hYRCNRFn85X18B602jpkxKka
nNU1becYF6Gr+WS5/XesEk04NgP0z5gjJwPfgfC3oeqQW6sm2E1gQ55P/xPbZK7/sRXy99h6u3ft
lkbPqnC7qsRwyWjKTb6iRMJ5LwAnFPeJq2V4VD8mNgvkprrUmF9LhKPUy1MwRyp8hB8XxByO7LbV
Sh61OEz8EWSXf3y17ZII94fTQWlas+YVqCasAcqKIDYgnIQvEvKITagC4l/7EaZCJMnrK7MVloHc
GNlKEssak8fe1NbeZ/BX0Y3ghG4japAeW3orDPiXG1WsMHRYGq9MdjTDsCUckrRDjII9o0Lu/6RL
MWpdlKWMVyiscS4R3KbJtZi2m5wvZqxGjS+M5nwyki9lEVebNq7LSND4D3q6OwADTAT89Qip/1Es
nY5PXeg4kiZ5wWG2RTdqKKDtygknVl/JDEUd9OaeO2JKv4YtN4ei6FjZ1FaVFrWbk6kjcgcyr5ON
MHL17q+RNcMs0x3fqWRwg7AjuVkgwTt2u+F9DBIhqPiWufeFbR7A4A6gdlHc3+GwodxpnGjt3Yg6
JA+esWrQJCM6mBBMr7nhMTbzYdrM/x0kNyRQ2Vls8wJbtfhUJG3x2jXOwD162kTN4YNjPg8B0YxB
xzgiaD8pdv5lxzhbiLdvoAh1iC+EILbxQS56TXMfsIrnFSgvR8V9D0D6WPKSRBaXrC5Xmv40Laob
sKfNJujTa91f0SjznfwCO09KtKgiNbg+zVOpqi0D9C+ujwI/VtYkD5TuHBIroF7i9t6zd/85Aufn
EvqJMp8r6ij/sxS1XiHOhRfvaHRtM1dAh6ki2PPXYA7+T6LYcYbgQtuinnkR1V6YcNlbJU10GbRE
Tq80Q0+ErbAD1DDORVV1nmucy4hUM5fBpdJKGobZBIDWLocjIhZ2WLWjpYIz0M/dLwn6Yo3V4/Ja
ZxZ1/ZqF14ZQNkkaLxxKb5N5uCphCL2dNsYhYMZQM66zx66sAfEnXlmF92QhCNPVt1bI5LTikEz1
ANd7wOkZPJkfbrKRKYY0urLkZzZFtw/EySgbsvmmVxgkLvEljIz1enIn4ZhpfqoR44+JDCxth6fN
IqOf/nx8COoMYYDojPELCpQys6bCEYGCYH0rm74UO3BJEEz5puymQzMxBQzIw7TMiZXQRlN+O9PW
Gyg7xIGFHMMLdR+PnDtADxHnX3fk55PwSm5uPdvTWmtS9HS3AODas3iXRzcTDE0HuOpO37FXVGtz
5drBlRGqoS5UNTxABzQZgjA06KE5AlgWu8ZvvUMRKcghit83XZCVRH+gT7ujEcVA7x/gsApOwNir
SHNv1j2qg7ABlDn1uzFD8ymKTD/D6qPahCY6D7WqJrreedcDFQ7HrfHjq81aVr6qgzmRRzS85N3j
68awFVR+zmZHcnFUV4GQOsgPdksPEbGDr4hxbiCsrFpy7/UVI8532lX5b11N9fcVGWPz45XkllF1
N6x586CCW849KICGKFr5qcYQyw2CRzHwo3lyLYflSQ/UzQgzTxC86kSKCj44DGwuhbNftDwTtnBq
1UeawFT+FdALhhUaig+S2/W74/44SHCI2asXqO0Brd0M27RClHFsOKfuUWWpAzquDgw/7GX8jFkv
Vn6OZAFymV63k83DuypB4PtMvcXAPa1PVeoQqlcNvuVUkb8+iOSQVck9CeJ7L90M3913K3Q1+UQD
CcxSRFTcw4PW7OUb3ZAtySIgHcDoZIOn3KOpOgCuoGKWaHHpBoozv7POrhGnnoo87ieOV5v4PrN9
+zf4yKD6TKyUOOYzpfzKcUrUtgsPtlhYl6ew6seUtaroZCNF3ti7gmpGUmNJxHZw2o2wBPkivhIq
/v13fKj+dfNvpwojV2K4QSZ94IHCGO0xz5C5K58cw/JjKq3lpiM+6mHpGHP9M8/z1uxIOc3JzAB5
YHS2FgnHkwbd9MIVLZPhQ2mS9fashW3TDJeHqF7IQK45mAINNAXuZe/pOGHIjRCQ+UEWJs76Thvx
sohrwTw6kiykuCku1Uf7ViB9xkrJnE8mrdwvPv8lsnRqR3oUCaLGyjOYt1meU0N1Lj6Qz58GE9bO
uHhIKb7ZJobRpSUNDHnKVTUCDqpnD+C99IcIIP2TeL/IdygeysCr7l5u3jGIlRgHXLY8ZLLDyqWS
OpV7oe0N3+5/EAh9YG+u17fHmqgQbKW1iRTzIwTlYDop2mIsVaVDu5wlAD08lmg7uWchyvnd44l1
+nlyRJjc2cqx7NMuEGGQgqr599tlqlPZDRAAMdhmWPiwTlrmlTSPa8AywziR7wp9debAwNLWyG7s
b8qWEYScdKKODNfehqHjlGvAIjVlQCNBK5p5Ap+OQA8jmwww2Vxsitig5IcaAIw9+OoyOWEKV83i
R2cpTKUd7PpyabPZ8tGKG2RuOOLo2nPT3rHwHgzp4eZpH6bQZzzN8qo1d5AImwJx5pKnUIfGRkc7
joCh5PFxoq2NyTdwD9/mwzXm8o34FY0xikCpEfxc1QX+Xz1x2sOMOzmVWrgkTh0nYwI9gPs+Irpc
1PQVYwRR+6YhU6/hWShWc7U8T0g1PMed/C30vHl4TfVKaJZMprT/pfdSu5yq9Iu1QJlJMhVsnJ4k
h4IW/0V1v1i4XD/QgeSOuX9mcODsShzt5UQdw0Iz+LOvWnY1jomAYIQdJ6UxDE13zBZOWzX/RWyO
IgmS0HWcYlTX1UqsPLR28Nya04lz58Jc+GcMh5mx+EVGedNB0ll5Z48b9p14uaVIlLC3hOafZh75
TIl8jkxsT44cCmHZ8qZX4+9hOBiQ5ym4Q38rvfCAMJw6Vmm1OzNIUO0Azke+seoAaJ2Hmjk9DBJ0
421XxsOUnSEGeFiJuJ5ujy5nTCyu4D4xAKPFVws1excyaDdul8k3WsD3wqvzZ22TapHJDDw14XPx
EyFeIe6Lr54fSiprmft2ThZvGD3pFM0PXpne1u4KB+4+ck1hvouqvTzXXxcSrK1D5cb5UsNvMwS5
CiV7jr4g9K85MCsRwTjQiGWoz+y2qkvizSXw4jzOi972vEPIUmVRjraaAdXQoygv566S7ZmwNzdn
eUU59OcJaIDVMyb6TLdfj4ZxGQshLVmoqko3jkRJ0r/eU3NuLafC3C/wceixW/rgCtX+vrftdMgu
oc+rTvNQlO5BvTIeN2KN6ynfKqVfocvfoVL/OLVcjFk+YCJsCZFHHyRlqUaWYKbiZ0MzDSh+AWjf
Pwglw09GFqPULyEn5CUqHE98T8it6BmN1cmX67+xt+h5dw7aEpQJtX6satQ6F6GsaoyPomFjKiRQ
+PRbSBXU+JYFPxQNulEVSWTKQ30BtNkIKNRfS3sqI2D7H6J8vk67dTc5FlevF5amJ2iCmNuXHevj
+vfUnSXjgi9E2GwpinTdJZmzNGVT9KIfOjDhaXQI6AbypwgQRLzaltu9Zwofvm6d+QTlaN3v9aFT
pEDYyd/zvZhBBwis5C3ORUQyslIsZEq+ktcd2DtDW1Yel6cx0qL3Lvn3nKnNJLpUUCTkcZU4zp6U
niQV2xjhLtbYvOqqhVGTXmjO3LjHqA1XGA3K3UNSENXU0gzcoWNSviN9INe0S/QsPLn/oYe7H+sw
XnK75G9WBruGwmpyp85y3paQQBU8loi+d2rDPKrCOaa9bvLImSJ4Zbn1W9GBnZE7Zr0KP1VoYFPL
H5C2rdm1nUQP4NyW7Li4EE+cUhM8Jx7roWgq7JItawLGQpk69FOWRswVfoEarBOmqqcdGZUlV0L9
azPKyxZ/+X4AUlR4N8JHlIVpt9JjnUz2m/TdWLv9Ds5z6WVipCQDI/upCKIGp6N38z03J4PTccJM
lREkWy5e8F0GnDOVGc0xdaOoILwZu/w8YgIxEtmybzcAKNmJ451fOCVbfmkj7SpQuxs8BedXkSoi
Mh0hkxMHw4pTtr9VEcNrw3+jFWhlPIS1sHOBHkp9oRYTThsj4OvvTcZNEQOjGEXW32OAdnE4rVD6
V+RvYnFPWdI40w7bAp29eG4siFwo4aA9MxQd7bU2qeSYO0I5kKggeCWgBSDNrFA0CZOD4V0WwpAz
DmIjPwTdv3rtLrzPkz4DErwXu++4AJwO/1CIyNVpYg+NVbM3DXOt9lgfXZ9R5xoL86VtLu3z5+/v
O/QcK/uPkWOBva63H4vHDz4F/ZhENV+kDCsz4FoAX2/6r/Kte0uoyoCgH7EbJtg0Zs9yrfDwQTFS
gLvJeJO3dQyOzYHbK5o8IdR2GLK8UQAs6dfdTCp2vTeOl4EeVndzUgqaKmKPIZLIJBd0GW2pJkJw
PDdoVzfZc+MVdK2FR0of3sH5pF67jiu8OxtBsFXbOrKdUoLHR6O4b3mpBUjtn2O9NghpJbMOj/YX
cg6v18XWBcQr2gZwX+Gt/9EpxSAYGG0ulS/v9PzCKP+pLinn0uweQidOoQIXTxEgHTX2idp0hrtA
LVR2Ao+W2juXN3nNLpxscllRJRUuwsbkHp7hhJ1zr1qLtSVWGO5QpqpJRo3byuis+Yz21NXr4who
0c9tKrXc1+tUi91211a4zOp0xa/fZF+2VbnHEwl85qJhztiN7Tg1N1GIz4gdKSM7X7evudy/7Ytw
9F8hA0s6/0tg2i/XE2hBJzopK9fYQLJSmirQec4HJbWAd7tlwRJNtK8w1IwmNKnE9H0eLrGWGsVV
3zqR23FPQfC4l7IzgosmVcuIPd16l5q2hMMwB/sK1oVvPe7ZaiUW46wCoCZEaARIfDiTHwrR4fHH
9BpbNN+jN0jqRkn1oun1micsXuhnb7LhMUTmDYJFB+S0r9pLKlFcm/dJn8nUKcCAmSJcbZ5Op+78
mp6srXYJK+aO+iK9gYAgzrQ4NZ5R2DMxhYkrGMVLqf4bU95nVkwhss9cf9y1Ir+lnbLSe4qmqjP6
iQgYKJ/dv6k4R7X4pQ1j9gLO+L/ijkY9WZk42Nl9uX3gIUfUX36b3H/mfDIkgbprdvWWJSEpWfPw
PwF0dj2K2Dl+Y1dccOVJDqFXCwJ5lXxtFFc5WD4S9qEPj314NJ1+Pif3rBiR3bnNJdBCvDuwlTbX
zJXZJXVBEXuqG0R65zvDRk4CwK4qZ8eTGoLoOEgU73HYvBQiom43EcNn3NS3zgLk73DfZsOvj2XS
5UqS9pfz0F1YKZ9UWM9zxFjdJEESiYPnLmI/Qec/Bu2zIdCKAkUTexJ3it++l6jvuDfwbhkFSQaE
vRsyhZM0j4oTld73D5g3FjfD0yN7j0yP5hxi1py/SWkyD54/3P3c6y3eVi7fx5DtkPoquuRMFfOX
RfrIvEcwzLjERAPOjrPQNGtMM30vWM2tXAbmdNG1eBNDkEwB7sxE3aSFB1oQJSCLrwh4cWH7RDny
CJH6WTGxsscMXIoChsW9YOoUskKaRq/KHRM6krX9sTT0UWi6qouZHRyKtiffqMo0usHTG5rGoz0b
vms2/xb1Et4qXf1K+pk79Zdy8CJBoOKf1iF2DzELnvht7tSyW4aaE4Bh63TMVipdj1XvXlixJWWO
cMxY9XNu46w5lIrP4N/QKlxOcDoxipchmj+x7/SKUYks6BLB7UXmdqb8evNi3UI3H9HK9IZGqAPz
mPCUJX+XTCmrfJJ8J6Bf8rZ5kCM72y6fz9o2nWCiL7ROVkVVIdroKojvxbw02SxslJzS45m/Q7hq
LDfhvgjhDkn+92oUZFVAXGXjsq7N5jsFOYRKSxHPILv2vfEv0b8hAwumJGuVjNKjyIj4yakekt7s
0ZV1idSECFCOWqlFhH42vEveN9QtS71aSBhDOm7P6ETz3UQaCPsM/9ad4iu3SXrr3ncurrT3CaRR
z9PYd95iE2rTIhs3L4Ypz6IZlh0zsu0MVmNbB4V9bAXm6GJjrkaurIChPulZo7p1wcSE/8YS1nAn
yjA1C8WE4YxrJA9U/OScUTUwVZ7VHExST7nneXdkHizsjPuKvvA1JB6HYyjG9GTIHZ+Q7fd9RW5R
Ee61tSiI9o5ZF0FSUbjKjUpcuS46kk6BbIdp2jw8DO0E6pGDH4UyKMwhxkJsgk87k/WUDCN89dN/
96nYMHywZt5OVs7zzQaoSYoMFOYNQfaAD6a5uBs8HavDKCHf6nifsb6yY8f5IVDDm2JI1s7aI8Of
4lfSASKBD+Hy/5EX5GXAJCZ6yYeJvPaYL87qTntBCLghBeAGTte9sI5z86TMqg3xqX9R8Rc/D9ud
mb4I5e0K+wiwHnaaidRo3FB47e9IocKa7FiYTo16PNjkzj64u1SOr5x8lasxLxssFgp6cr+/X6El
ddMM6v+MUEtlAGRYT0092aTfYHXOzFq3moLmbxhEdeN5J6jbxpHLmSZk3BuSrwWjQfSr2VBIGL4O
sROYpErcUTUtYqMsCL6UdJVXixZJfNpGsGm4dasc5nx7eOpCpqoH/TCtsDKmVCfaFGczdHvOkw4T
hJcLIGu6vVC3BySlXRrlNDG/YpkEqJc3l+qhK8XKatE4UGlbCizry2il5YkM0eLRLNBlScqqCKHK
bFfRRVI9HI/AYCMuJco9V2unhe1nLNjkEbvbmwU9QbxJNl0D8kjxydDtReHZgYsx6NQdgsOeN4DA
ckQdrY4dBc8Tn6L1W8eTT+NEYKtssnOWY4lMIgR1sQTWwXNyH9swmvXh0I1ezlbzzq9nwG+atfB0
2sZdoiIEZm430URFRCvcVrVCp6XrbglkQafmH3fPqQ/3nhFcjnQfTU3iqkBks22ccvUhbPBT179S
o1cwK1Bgn3+WmX+ChvOgxnrExlVm6mBu8Xf+xEn0fEaIT2wl6Gv8C/kcuYCDw3JlU/Hk2mFr9WQ8
6wcg2orkq0iELft7pdJf7W58yHhOrIdN6OmK+Ob1PmnQ01fggm2b3+Vt9pwtpRpqmhyM/fqg0JAP
9drkEqbrhtgcudKjSR5ZcwQ1qJwsnxCRgacezcmJzqjB7czcLp7UMfb4jp1R60ibkbD1v6exSLue
fy7B2/ApHxKB0Egpp1zlmSGTNXGyA6abK6at195Yp9MIovWKpWYM/EDsmLqB9pJDmv8ya5NSgmBm
xQHNVq9/na6cRw8BF/uqmJYnoI5UwtAfmkiBr4sAYdWwMUMB/oFg4iyS58RUfPPNM0wAmFi9JQ3u
eYa4ZN+/KcB22D97ZEdDJH+hS6lF7CXZVYVUs3PLKUfGPaCpT/wSRuN9mGgudR6LpbP3YEpbs8Sf
gHaNlSMVxu4UcmlkMqvqL5v1LQzBljv2DEP0093t7UWJ3ujQJvfY4SaGJJ0fVZoUubd7oiVE+E0e
WhuG92JFKAyOz8ANK+X64FORWTpcA4J8kH9y67slnVl5aoF5S1eczKWGEeybANP9RrY1CHi+Kt7d
1KUl68SHbtob2TmQ8EH0dVZ1fy6i4oevZ8HTmuNN3loSlpFyODTZAdBickrKDMCJmAcAhwuTiMwb
QNFeCz2pTY1CS28VfTHFUIvK58pPq0R4S6jgSGEytIrz/OWppVTMMDgondH78jGUKW/upjxXFD7H
dJSPm8hBcWcTNQURrwqrakIe2dWKqlf49FgorsPvUIDhFTrMdP4MRwC5Pi2+utQ4DQyfvq7Xew8n
GLn4j3RUpzvfJRnDx1WopA4BlwAJH2QY+Xqye/vXR4KTNJQbf9k42CGm7TFt4FtmPVt2GjMsykmN
0Q748vPnI3ePzF2/z7O8RNgRi8tAEd9cKnuT9qvRkLT2kzJB+qb1SoiFdWOIHtYcE3uckE5Avd1j
WnCrxfzcHjSBcH1FehsHBQTBQLDSB180lV6FFcgqJwMvuv6ycnh+Dt4pfxoGt6Lq7TD0iybSKQs2
gthTeKKQASGjMtqANnbsozXJ7Fm+SAklnwVyhyMZ1LXdEcT6fxZU3ZC0msVkjHWBJx4P0mWA3lzI
QJ5RFTrD7qFlN6rV7HGKK6ipjD4DXpuIUET2OcjUl8eNuhqKQqZBglh05WKg/sVVWT25LJ8XWprV
tjVs+LMAivdphR0LODFfvcLQRriD7QdHUtKkGYGHdgNjIR+hg2N/Nuk7wrXNbt/i+j3MNJ+O1LuS
O1GcK6DFOVXV22qzLyh7ycUbxoM9H4lCikqsxRbqtqeGS+MU+tkvfNty/wP2qasWN2gz93R5JWnH
ZrUFw81zCcLyIMEbUvKO5HjDoqiI3MU5rLbSqFda9gh0cyVO+skx6ObnytWuh5/5tQBmycLAwLop
tl2XBQRUORod/A4WmNH3HGYkBw0Ba7ZYHNXJ7K6LjJWQdOz4krdcvcCltig9mrM1kNFlUGWT7SEh
Y77JioUPGFQrVh4owU3iOM6YUnb3oyaOeyPAQgmFzyQcvyqsB8gWOTqsfJNafvN9VRtbHwIluM3q
06PzjWVsClqmUF6znFaSKpqql1hCwzt2jpttKwIiPwrqHTlS2bFfXwS9idajq9FwWsC9IEfzVuWf
8x1kwVLlaTi3L4wtkZAHAOvhp+psqCmOOasXTWG5l/V8jigpu6OKgxWxdheoueCqV1N7EBRZQHcQ
63TgzDRM2G3ZJg42a15FfqVX5GmCls7Bf9OR+06cBrOv4ZBU4t02qDWVdR8DLo0dOsuzyAgzdMVJ
cq1qw3Zk1Q0TmyFMUXguQ4iJm0jOJ2cD2AV4Rxl48Qpsp9gXxD08Ve8HEZIQRW9x33aY56HAXwIz
FK6GuLCjZOqGswt0SvdjcTnA7NR2r6G6l2WznoUKbCgyP+hRE+glA5eIC7hxycuI0VbClqsBuF05
Zy/cT3gTXJS3L+k0Ecptv6Ht8qdkZaT1b0RELUUZSoAQCmoPMIxPcvIaKaOmc118QCfcYNJMagrj
ufnuCyDu0f8I/yg0aQkhJoF8LhZ+ExQby+giTe6KPJk49D6EOFO0vpVUC+ez0Vw9UG89BMWL/Nuf
SDVXqhgmxV3OEG39ZBTOYnKV/WIfgIOnsREEYc1vEDHP+3tOw/0Tq9Cz8P3nY4Ez5jlH3xar7an+
eiKCWZE70VccBw5F45wj7P2H2aI95BuSUILAFuhXpWCqUEVuBcqV77VgsZ/LukjjSe+JJhHPGljV
YQW/7vznvaDUd/wYfgguF2JVFwlbkGU4aqbYD0Omz/FF+nBoxODLOhki/fDp4KeYqS4pHRUM6U3v
hT4rw8vNV3V5lqMvnmAbO7ni/Xf9u7r4OXZX+JOfGFtx+oF2IDfkomdjcTPTuY6Y/uU/ZbXAxdgh
ZIboM0tZICPL6oZyNktbBfhygU9eyrK2zyQJKh+cvED+bG2UWS0qpV49L/gxK3oSqI4dc4VdxXSx
1cevAA3pw798foX3uTixtSFrZcnSQ73dLCphvWfQITCUbqwxrza1ZS1sWblRZvJwIk+xVZmgc1oQ
L3nna7lXKGEl4lZrmjpEtnTSFcpTqpPjW1eapfiEcEyM7HHGnj2fOqytF+zzvJTXor46gzd5thr3
sHWXSOqoPaGx743rmV9gIN9w8+26YOZEAwgaJCDu+u/YllXDvkAicK3QOXJJLHMancFJOQ6r0jai
zHyGHjb4++kQRaMcFlZgM4Vx2ktiCReNkElmCmn+G76TknkvMNLKr6H2tA0BuWc+w0DH5JwwouhQ
S982sawOYO555Ki1Ys703IdJQi0tIlFq9c1Q5+Fl8TPSCJ4YOqEgtj0skkFUs5GUekLx98NnBm0z
NixIQ1JfVarD3/pTcWfSZBbNmIX0bhNdptorlsxzZjuvD/lG4qaOtZ20C93/nVD2ytNN5lBKGQVC
x4HqbqcHd72l8OCcMklls/1RPE/zLJVlIwPLZhyAh1PxE9JTKlW5oM8kHqS0i9oGECS6+hoBwa6f
Fve5E2CbxpkIZbx/4tBR0eAlAb9nqtXxGEHK65Py+m4iL7JU7q22LgBviKYkEpHLnbaxRXNVQ+DR
IQF/Sc2Jrrc6cnqgCmkTETDIw5TqnkDjNMrhuCTxDdcxCIlpK8RBgZAShRVA6YC9ivAQsqK1a3/c
Jrz5F0e8V+Hz388c2BFap5KPkEP949pwtSkIqDAQfwdYbPwCOp0tjc1JYPx1qk/q+mn9n/BTjg8d
/1JJFLXHtITO1VaQ50YwP6N7qJ2HM0VkrAvmgXzmbPJdmKXg/mO2zUb4dTpLVySfq9Gu5vP6cH0/
8p/esvz+AilajmlZnhpSvqeYSQfgjp1KEGTPCUnkcyZkTwb1GVqO93lZQBl8JVTePKKy8WJ3Kjn0
1fZ+kTqBPQ3t/rPPaltW3DNf4NW9+G5pv9KUcQUda7T/L0hq2Mfrr/r7jckm1avtqfCzfaryYo+s
4moJWEiwRU+w3GvXgPc8fVlC+RcOKySRlM+V+7gkXMPG+AmjOC+mGQuxCo6WCkRxJRs3tpNO05VU
9UCKzbeAouVN+bBfVUA/BfO9QLXAmXv95QEUhwmLFquASwaKlYV/9SbcR7zzJy2dXPXsrin34dFN
2bSJEoX3R2QohQR6c+V2tNXt0hROyxC93JmU5Amu/c+oxXMKzSQNKdD44mKPZusa092zX6zypCKL
zYhh9H0/hG6IDeoad5PIt2NNp9CCRUaN/KfqB0TlVoIxdO/6jvuDLoccXOV3SJgbY9twV7HQ2BMe
iCNjjGfaSyMzvrWz5CcAecE0wsFlGhWqRiyFmnCgP8SbdPi+kAEiTLMNmJuN5oeEVmeGcvGooC3E
Furf3TlMAcxXA/UyLy/zxTDtU1oBJ8JYEdAwTGsDGznn3i3hGIe06OwTx08IilUJH/8T0/1Gg7Wc
eft2UidNob101XBW9hoOa7+lTNPvJ/fmP1R/zFkDOKe0e5b9XX5fW2YH2fZMcEqU/5yU0eyEW6ww
K8PcEwI3EKdShZZKbJjGOks14cdMv3MayDIAqFk7VP0bW/Ehfliozvh2Q1I3oFXnb7/Skd6aEdvl
HWnN3+kRc+O1hz6qYW83KsNnWLZljMkIUw8R12FC7HOobGuJhwlWFuaMVwFW0CAPdHdadAf+NpNG
43JCOgiMDTXca+LIY+RQZYIYJpGqwpPAw18SBo1j7Svh2mnfoSfjdU2lLUE75NAbTY1atab74WJt
Jwljf+ZPafCCe1PQn9NJ1Mq57FKlkJAJ90z21okEDFmlBxDzO7RaQM1cKsJzZQ9n1VhlazBxwQzh
wOSkl57AAxY1wB0lsqZb8FQvBin5Jb0/JkzLaqT0IEojoR7ywg9p545hK3Ai0zJGe0jm3LN34q0z
X3g9wMfFBH4ppb/QScAAy3HZJzGbAAg48xHcjyRLcDJ7zZBLJ4jSsVB/r7FxxEZGzfSHiE30Xrkz
urSOMJaxowf2N3BHI5uKyXNSZzX+zETfi0AoX4qVuk9vr/w25N8tFp7ggqQIs+zeI0kE8IxZ0+66
05XHpM4tslRM570yUK+PqaSy5L2mAzjBCNOJc8eFGT0Et5ltDNtDQm2BtaO4r+R0HQtZktgekoKX
01Nx72WVS5Yi4AZ4pPYmf6VYj94rJyh11GElIPEL/7hytNG2V7kmKv6zqy3kc6A7sm5BJC5kV6Iu
w3mXe/Cae+nVCM8nmlyWC60t/IBqYgbOdV/9VUHM/u3U/E/sdY4iSqBJXvsA38bIQCHGov05JMgY
B1bunH8tNtx1Y1VEU+emiqFXW4Y/jHEIJ8RYTNIqLs4u2PlgE0GsaxPMX+VzFFR3cOex6pNDT12X
38gKkAu9D5EgHigEWqpBUW4fcF28n5wFLzC7NgyF3kt6qwCSekkAkJRHgog+o8HC5J6+/YBNpC0A
I9dYV8VfYabUJvmiJPGfpEJDjzz1QGIRe8J6B0eu7+2uleXC1/wP1fhcOp/5zJ0+yFZhtHm+h/XS
Qb122m2K/tk599zNo7/itJ05VU8xpF2wqeXqodLJJdC2K841FpPRNSpivbspdXgEPda2a1R1J4Yr
IoryM9+Hjt2EXh9qWlFsqURgDUGwuYGlHhrL1iQwrmVnL5TRrzhwhfOxGEmpYM2dNFR3PgfuHYuC
3MtYnvE/3hzhQ8hWaQ0YHcVpae3iKT18E0ZvLnqLJVVybMqX+hXxjWmpwRXViSZm+AS5O2VlbHOB
SbKAHlxGFJhB0c5Y6uB1PxkzaJZtP+q5B4J2KDJWV+93jjxEGGcBCxD/djt30/Lp3FY8MADWhBut
EoOj6LzIsDQEfFupuwnj/WUE1vLXzn2ErtLO3crCK7u7Lk4kI8byh8Ynsv7ZFMHtmlDQ8DMLMbMo
IK0GXxH566PiDL/X2Zzc6Wukjba7G/Yb23gsqaL/qt1KbKZoVUAD0531NOcvLs78A1QnFaBuKWIv
dFMeZgz5oNJ1gbzZcPxY54pB9WBASaFCTWNAuj3OP11ZfF4hONoZPi6QExPFbLy0PPX3wO67t9fd
qPfFqkF0wZ9BIHIzsXcqLf0V1X/xUxPTzheboNw+qdzI+V+Mut+TBzHNkEcKdAu/E4QLjiHM3pCl
qVz2j4yS27qryql0VoCYNt0vkH0tyGHcHqfGOe4TJoIrAgrNOB6lwEa9ZG/AG+gu853YPSp/oAlq
njc6WrQ2JkNfFQ+tTxHoZ+LoQln6KHV40922+SmX01iS5iImyZcDxJqqwTSc2zR6u3NdKWlDbQaJ
vNGLZweyNT2Tq2Ao9pGc6/I2/TzOB85DvPDJuEqj2+bxNkikbLD8v1aVxzm4k7aV6o99wUKmMmvp
pCORIXwCAf0hCess1hSct7JN7LY1/5iQhAla7112IM6zmGZ4NUY+i7wMvcyX28PbnTBwUeuj0SGa
br8NBKaFI5h/DpDD1wnNVkyfh5u9X1Rc4BDVed4wZ6CgudGQXMDwO6IvtUyuVIQm1VIf/8I3j8TQ
pFXh+9OJxGO8FjeLqOHEO7NS5VqKMjM80F7Cz/HzqtBr+vheLHtNR7Je37g1HHNocUuDYHv+IIu3
ekiO+ZzUkEzp+MM5NuQnkM39CZdzaEuw2e8Rr3LG2tVQNHvWyo7tZ97mnhvmDdu7sjEdlmtkbTA0
89ZIWLM8AyF/dlnA9P0Ix7tXFcKKvoz4taUSzghyl8l/2s0dN0fjsRd/lIO548RA/v8qHwCihN1m
1+UuBnI3XRfqSvN0j5IxAy9CHRj2bvBRX6iOL5oQmdKsODsoZ3fMb/or6FE81WkcR/V7ez10QZaS
LCm07YnPnX4qLGUqIOpFKC8myADxm2zOigUyFPL0t3dMmm8NabucaK70ND99gFb6iQuXA2A+6T5H
zdWaxQU8R99LSYguMcUWq8g6afbpJDUO3Ps90QTPN0TORDC4hAubnYFDX3F5H/huWmf+2ZRhCqKO
bPBmjT/4OuAOeHObD6WmDbKGMMerNZWNZ9fOU36OsHTKbvI9HAu9F1F5I8dQQHblomOOY/RFdtgi
wwFciz1mqelPRSSFanIWZgwvwePnj8Ucw3wLmANxNs0t0psJMbTNA1Oyk6bsAiVOUACq5/60aqyq
8FaGmNVox+gOfR57L3HOI1nAelOcQtmJWWslOCPT9lJ7DB0acG8mIGNU0YNxbr8xdrIWKJTVqaL6
g/mNrMOlRoYatYrtCvTxf2cjQCsEkeGvc4C9rvQXosJkl+q3pI6dpnHZpG+RZOHUusfJlBpavkCg
FRwQ/BYmQIjG7B6WbAJ8TRYpXFcFG1bYuxPH668Cj0WmMHKCSiphsRRe7b8Qx4W6JpMNhqtlduJo
EdEfO0JLs6UtXjbTLkDSjZG5TPGp0lQjtMAUOcTYnhNILZ89Q+0cg7E8SEk2AaLOV/zjYPbsAbyo
aYBJ72i3pjx1ysYUYc6h2Y1XGdzYr+x4Az25hJvLDMzFQsg/g3TbMpTYHAI2albsWtMcqKjO8mfL
Pu1FPwfafJWHpvySTdt7QSGwiYVF1ceWzu1jgzL2v/m4mW3582wyn8zh+FM63k0Q2e0bEjr47/su
HkRfUI7DLjIYqClrpBtKnaCeBMjVwJMUNdb4DhG2pxHSQevC+W/WNXFdyWijZdnyDiq/yJrYW6v0
0yldicjFdLTkbs01x/4IHFX5J+tAsy5H/quxvtURi/Fl38aSE4hOysqzDYygZDkfErF9TxzZvin5
kS1NLdorPwDvHo2Oy1WS/uHAS7CnvnaSOh3nEfh3dXQJy6fLTYKP9wyTI+L7ySguBrBeJ2RaqyDf
EtXA4qa6yqpN0ncM/dbRoDn99HMkpTbqWVgBFvB0RAtZznQhu+zN4akePh2qpl0fW12izccFPhkt
RaB9kXJXMC41dnu/AQ3Q2psMduxU+F99LNHglfludMbCSAzNJ+kw84mqmDQv43QzSzqcy8q/Kk+K
1WcpSJ19lMBj/I/xZZk9EkUiXaa0T0wkbG794sm5DbgQxz1gXr4vkdFsJawuAl4MrxhBhMobrzNK
fn5KWLryfmqZvWkin3un39b9KJnnSTu9iNBUoDpEOy9iAbtb/y3dwRQ8v6QmYNjvpImwE468/rdT
kegOSbznZxUsm92bAiLY2myYwAj5c6gx35b5cckmY/PAFAzLtDPJ3aGYxXpaUb0/5Ci7IqOny9a/
eXrB3Hyz+BO+kdip0BKptaxGu1im+Ea4mjPcBOPuHSGo0hXytU/rBg+5dvTF4kqHaJYnjrViHgpP
155G7hCgL9rZuksAkI4miI1jEzZ/SnDx+3OsFcQFyim6wpjJNnMTzlosfKDOtSJrq9KxjPTfjT5m
XcNtUPBXKzh8OjWhgW567B3YT4TGgSYgRocjH/8KY0wjXpG+RMkQVSOXPFdeL4XnAK6yD96VaN/b
ChRbtKWaknxdJk23fCCpxCEEe112UPRuilhgosTO0Wspo+sFW6S0aybtFSpumDzvSg2Dqndr6K2/
V7YgQexmr5hHoYv/qIoQDP52GscNT/xQm9TVsFKwvtr1lkJxBHesvQT8SmIlyX/3wHjWRreOi3Kj
LZOHssXm8/dbeb6llc3+tyFjHs2Cc5fcOi+8kpT6ABGOZYIMrJxP6TPR/H/7B/dprGtNkJXwWHBi
1QS9Ao/UkxwxDCU2HFe1hYLEC3MXY482Z/ahSEEOK3bk5LQZlFsH3hfE2WE/MQO6s9hZgFpJN5mp
j1+hbo3IIScayQzII+9L3sOLjlBqFJDYM97XiMhqM8/ZtsfaoOfW6ndYcnRvBA9sZTMqIwGK+gUl
63HWA724EVXBKfzUDaBDxLJ3MtR9K1qHmk8VqGuquj4br8zmNTNLwrh8L85vxhAqNCh1nPyDoHy0
I3qcAOVlUXs8takWzAeLlGzv+oSNV750mnG8w59DlOmmQw2BnoVL7+pd/2WxLtzta9ovmPU3eMi4
qCsNnI25alJtlPgMdruZgBaEvpQJWTTgVvOWncbtoq9LlkM2M+0TIUxQ5EP/QGA5e0UviCud2fPQ
GZkvDU+y1ZkTAq7bLRGbiqHybE82PvcSw7CAC6TmKfeFj1qqxa6k6EcxapxMen3ORiK0mcpW7vAV
32oK1YsfC6LIsUBZd/jN4TdcnvIb+xeIBck2s2sq2vS9khssCC3CV+z0hY31l/GPdECJOihTGlY5
7O0I+NzX6AzvSqFc+6fSszzImW/GZ4cmo1b90ZMi3co+5mTsR2mknV5WgoleaVpu8abDfVONfipk
VcggbUDBnXTjGrlXQza9Eimf8mSlfrKSyotFsS93Rgi4q8hlspAB0EHgXqG0Zg9VYye1s2N6/NsY
zpz9lYR9SG7hg/wyo04+0xN2oqR8riF5h1CF5xeR+F3PBNsP40fuVy450y0srMlyzn4t3lT/Vaak
UGytUN5Fd7nKZzQqK9Yk95YMTZ4CVAR7qD+jgyNFuilBCnG4Nv6A8bzfuXmapkzkDa5kg+0Vdx5d
9OZe/UHbKgNOkRTHKYBM0sSRj0+nKNqirZZPyW82PSLcG/RXGCGeULw/1XO1ZVQ0hVzwd8STFe+P
CPcn2YfqjsS/bD//KImJxdeP8vcf/JqRXsBa0xEVfRhfw8Ak5l7AhwBWcAfiz06aIZuzi82BQ6XS
hpxR8Zct/TZsiSvdWSZQMnfxCSgaOkulguSbIYOo7D8ze1GfRhDeqHzexvTaJnPts+RJ8gCsQUui
+qn2DJDpvyia8XICZ54Rp1fWYjNkK5vdK/iR/rb6LioKyomjybFVPP8q2dRiBg3ZzwG2DSO9SdlG
WrLaU5ixfQu6c/0y0VMwXu3AOWYHD4jE6FbhbRtoDZcNni9Ac2bNmAOpns9pLg1vtlgbQKqmwam2
NF4BSxBH28zqQqdz6XuE6Ts9J32bet5pAKgasAJ7azDjKi5pmsGTaSS1XOplU1C1XNUEjYvCQnCt
9Ym0ZgxGzQWgX+8UQkGTh2pIv7RztBuebQKUmG873Pqyn7/BxafGi1kQiknCdZvFHHwQt/J/vXy0
o1iDXtr0pgwHkq3MetDILqVgGgcfA4raauwG0Mbdf9BU4f5apA/MpRmc7t0nBvn12heUHCBAn7Yt
sFgZ0KyMWkopKe+VWVjoOgDnBtLdldlUhMDZvTyRv9lkwxMHntzX//6TK3C5Y4s6EHSXtjxq3Tj0
HJTu0UXru10MDX7JR1TPLcmICQlmRUzJmC5Dv4A2HSAykcooMyKfdJyn8snFEppNAy1tHT5sSE28
Pp5UgpgZyuHw704YAkHs99iCwjg4fTctiJqUBG+YyE5j04ClzD/5N23idwX+L5GjCo75liCsl7qj
H8OEdL+S+ad9iBSbvd7SdHLiSSCA9ZtsfTRislr/3yIoPzUe1m1yYwrZOaWJEHUWGhhZq1TZMWMp
s70av7kjeKUDa1FXcyMhlC9sk53DXR3ommIZ8MNN686Yc/qioULZtBfEKm1lXREfS8kodHkJDrvR
uEoM+Yc8eQeiEzTyLf1Ne8qlehAIByBDMGCQAMbzpzvT2g8GX4s5xwGS3ZBVUaSO5DxIHa0KNqF7
bL5FzfYr/uIIKibWfmXepxb3r7yKdQ+4ezJtpypJIMOmT9yHUiBBJSlg7AKP8fYwn2HiT9RJnnQX
nTnpPRNiJa4tUa/HfLeFGhTDr6yDAm73arJjyG3wmdlU6/a9pdmw25NijYiRvNu0eQnoKlMZeDnP
GTgGg7SMlEgcEPyM4d1e+PTva/MXYJoL4AwTw3U3UWyX47h3utJ+k9AV/LFvfmhfH5FcWfwdN6Cr
XFW6xBdoGaaIoenP+VfyrGT0wmTRaFn79/iulU6hlMi13s5RaO3yRS1VxuzEQkLKw2km3X8NQ3YY
OAZwFAWYZu9JfCM2Yiw2iu3PlztgRP27+yzUj2Yxh8IRDp5OSDwJ9vUkbnKVsZ/s5QfgBuAJK9LQ
F0/Vv/i9vVJenPkXRQbyN+lyiv3xfTCGrqzKLX7I5SbWFmZspALP9t30yDTEQhOEpqAwPvmmoFHm
1DW/5FwE5J9WUE1Ue13HZh9HZTSHZ0Reo00ACipV1Txtc37rp62pc3PVlpSu1c0F/vpcogJiD1ma
HWpeE4Er7Dwjq/jDqvFm0rGZZiE3kiPOjwpnJ2AUt7r/BTg00N23lkXKTUEherJI1Vy81HbreNnX
uT3kACwhDeblo1pobs9ZjgCAtPwEmUsx68F8NudmsVlC2yABK+27k2pPXDDJRBDvLyJnLr78HIQW
87Kp3nUsyz4mnnVEkzpDLP5WDpf6ZjaCeNsp5GV2C+nU4A4BI5b4KVPT17ZZr+lqM+ZfaZlmjFLm
3eG6hz93tXCg/utHRoDlcH0LNFHgLb5fe3Cyk05czgsATW9jTSIX4vG2LOgS0ERmdgpAJIm3xFFu
G0Vv+oSPmcbOTgiRWTuKMzyZUp2CUR5Psrsm38f57gwY9vhCWoL2JzC1hsCqG+2tsv8p986hNuob
vmWw6YF+aspwOAW5Ct0SD0bFCmvKQIJZnqlC/GwzfAyCwjrerPwkUJQAgLcw4JK7f70eWNGbdU08
900ZgJAPTcfZZLIbfpSiR8PNIwzHH6Ssf0Hf9zUIo/Pv8rSr5Y4E+4dyfplay2z+ESTtaOORt0yf
yWg7XCLsOEpFatr5xLlk7BnsedD+/YkVAgESYiESAjB/86pfCBm765cvaCVuuxgOYnRKyMqEWwks
tr6ogRow4OYYOcMGH90WvkuCGgtGlfEiynSXMNeMcmef+AgzrHSWU805+CYogXWwvcVW4w0z834w
1+5Hi82LmDslqkb7wWJpT+hxPrAhFSrG1EafaIlI6L3HpEs+d8W6r6TIWz14wRBoeX2dTZO6DT/s
VTsN5bA0o/I7iBbCZKl5stcIy4KeeZ9U8OXKkIAwouujD0Q85dEan92oo/qZRJkVKxaodrjEuAwQ
Dchhe0P0UFM/6JVOjD3i/sLpdN5ZWCWbm06ALmEL0OPS98dztuJ5YL5ddnoYOAWN5VbixdZtpF6K
CIktrDaF/XRaot8Y/dvJXR+whMEnUDSC25i5YiresMN3va5AULig0iQKj9E0STL5FuEOnNgaY1dt
/xO3IB9Q94N0O0vbD4XUrmbAYwliNZc2Aibh7S7bgpKgPkf0r0AkjWanOU9UnOICNvAb6Mc2vnF9
LQxikg1IfN0f7GoZ4QenlOFZnm3g8fQv+M6A67aJ+6WujBSf251eQN1MEZ1QadEwPAlvlOQV11uQ
cYD4pW9PutND5KNHf1RVKSh78QgH5eHDukVIDrA7mt3RmAw0WQpMU+ar4fwvSle+5s906dONhOK4
PdOZcrudDt5w0ZhHy2KN2l37ipf6RV8DMe9V1tqS8jiMn7U4d/C3aCPnriT5M7OPd/0peiRqgTRB
t2T9SPD5kPYGMCaf3SAk5rs/8hluhmF1QYPEm87lh7A/uvRuTL7IYo+gUz5Uhm4bmbOyC9XHzQWo
ln+84ig8it/87/oVdLYTOjgOqbtQlXUIXnx+6EwmRThpcU9eVcTOd8TkFQACl5K1TDFC5aYBvbQZ
G/REUlcJN6zbSfxd8yirPJ5vq9rUrNbz/2NAgCGbFEo/ls2kYQmrr/NdXPn5ByOER7JoqeVrL7Go
C8gQgmIYlX5v1UKeYcAMWJd5grJ/sqPdRoK8+pG1b7I3BaV0sl0u6WplT1K8wtVcPTDlQZak3VdE
oa0b76gsIZuT94Apljfg6l42alcbWsLUdccd1IWn4VEWEJx/D8sAjTdCQ4CRCBK+d9v7tvVfq8fX
0z+d6/loARqXWFPwarzvUWGgj8UhhqndJdZ4yXwlIeDXksXhTmLR6prolmK5uCPchhFdJQB0CdvT
k4EacqoXgIpJ9FDK4xpUq5LcjU5I+uGNtc1eINVvXDCKIkdc+C99W+5Sp4XmTS5izLLe4kiKR7ef
ycUcuImbnUuJOOKDue1bJ0Vz78G8SwNXGBBRiWN0ocPRWH2kEFjeHD+/E+1PYBv/kEahUHh0D8CB
2+ZMDzyzHfilEoO17r4R2hvMF1TmN9KgZzp70NqjVUvu1sZDw6JC33/+ERdbccb05rGc/VwAAbNa
kVg9awlGNmWtxUOLggU9lCzP47yNWuNkvYDm+hOj24l0T/UhAY/iehA7Dk6rPTodxyG8lERDnFm+
64sBgFCU+jIkJdsRtxHwmS1w4tbcVmUZCrwJ32O/rkiNcKCjFEBqTynpxURbumQx/YQJ31tNiFeO
WC3/jZq+0sa7Pf6L6NggARP7IQTm5OBnD5ksz/pKhuMndsMRPV/SD7hILY2EJvTrXMn5Dn/Fx5u3
gW+JNB19vsijPC+biLtxw7J3u7iRgceVAJOXgG6TJIQATl0YUZPlh1XrPsKPLKKdno/srGvZOWqy
TgQair+0hgBDFyA/HErMRR22Sx0iNeLIQjs10KBWOTzGedzZsK3gY8hNPhydVkrsy1UgKnJQl0GJ
gz040fKCUrtITR8Pv2mrO1XyLAT3X8/8NOwgCcXDpTy3jsKr7IOTjUI1yAYdCBQqFxX/onAw543B
EBwGzqnXgHFe6T82yo4gUBoUvhQ+pOW4NnoUJWkicQneaC22S0rw+bhFjpbEfl2tT6RFFACphas9
SYPfvZxpTkjzqI28bx4PxL2Aj1F7n/dNaFFN2d1AYbYxQqvnqze5o9HbQD2Jg7DOXvO5Co5M+/cz
L1I/k8XVMj+/9bzXKqTiIKqegVklzG10VEEfOqQWk691GhwpXdNub2wwLWWlSmX3CCc4B0K3Mp0n
K3xwrVS+BwW703QLQ5EQxqpM2AxI0/B7xxypO7iQS4vWA7+baiDD7Ch0qWeFjykEmKq3IG4DHkGs
Wv7NoA3jUuOumOmn+ch7r04vZn5nHp6MNENIbtkzZ150HdRBog16qHD2VnNxqnxfTkmfTF5m+ddw
3qiL222bsZQNeop29OOxRsMRIpe/yHcCKtuBKfW7tcmknZjmL9EuA6OSLzg3ZgsdO0d/1U8lseVg
WlAcVxup4WOrywFMqrtQOHJpinRIUY+BX1QTsxcSTihzEVj6D9cu+WfRyd318GcViKnIvjnzc3AF
yP7QxUwhvAAA52h8DHQnDs5Zw8LrXuq0xIwpmbL8x+ztEZYpv4tN+a8TDtK/nn7a9qhjihHHGJM8
VtMOl4HLks9m8qIf8dFAd8wAWRNlnbilSVPdcq3leuRHnQKM3XszpgZuXI6BE70UB2fyI1xauh2a
JWY/c2BE673AKRGcgDTvULLOLTD0Dc8EF6iW4bXAiLVkdfKKzTgC2rcpCJrBJGELWsNxFLwl62HX
/bNBAUrx+kfcGsCx4YQWIVWlRgsrW8rBmPKlssjN7sf0EUr4Tf3gI4YUjIANudJXMQcxukYuGZNB
/6hgpW/OEhM9jx723YDr/lH/ZS4NBpFWYdUg6WEBCt9fk5NXnhPNm2bp0GvRekR6pFdoO4mWgnZ0
qEaKb6rJoGvHaYt0wzXbTubcLrQVvny3ZZHYM3L0gffKPoX3VcvBVSWpDtWXmzDE9dznLgH7y7yb
exbty1Cd64jg0/0FRdIcWEa1O17Jil92oX11Cs7aVDGdYUtVHPs2yyEylrOnGB1e1TlSmqnJq4dc
4Vs8TxFNeVnR6iwBmWk3Nvc9Xoj6EUZ+QaNUVu5ccvrqm2BBPbu2uDD06s+tYchLdZHnRutbqtCW
dUJtjUCdEOyhUkycN9WIUxldvqn//XxvgJ7XAKl/uMNtPZans2OgGuP2880X07iIZKA9bNhmPbN9
p3nJo5uKv1kPqUF8zfjEeI1vJypJAcVE1b7XdIOHsn2YwLUu3hJQ3xTJbRIcC1RvYpEPuehWhnsn
VObZVOCovOoCrQMItNj9BPXx6twnnyjePheQMmjYkqLCwHdFWb4U9UgS52wD/rznV6OIrH6JDXU4
q+hqG0GsrGp/Naqe3OTZJr6S772O9wCaBvGBqLp01FRezMLlLvsibr73emFKYOGQdciFiIwSbKtm
WJJHVr1sMnTsZKCvTBAYMVLFaSqW2u/0s9cTMXF1uvT4HdXgTA8A+4g7WcuwfBzoOpTrRi2m+HsZ
4yNi2tPTk3Q9tbaJ15PQiG4xI50f5MQ6UCJ5z48Pclzr7ssqiaQgM2K8HjClstIrs364NAvUpyc/
CDNUD2T2NsyhX9GQULJ3Qv4oHFRb+KovZ9jj4nBzM3ZeOpY7FhVgTfrdT09yWXlku714tDZz7WGe
0R3HlfDejzGC3glg5k4S4llg1Cu/K+h5Liv1chLg6bd75YwhF907/o8D2zR1q5v2cvHwmHYxrJlb
T1+csqk6zYHkHPPBLmCO2sTO9LE+GZuBFQwbmVJQrKfagYyVUc56erCQFOLzIO5Hm4E/j7oRfDr5
YVW/RxwQU1q+iDCEKqg/V1aJhJ9JsG9llnIngqvR0nLzNuRHEpWatLRfsTCa0zh5CP035BE/Wg2C
SdeDKUK2o2KVI2nEZRQFgnDEEcnmsgXRIxF6Rj3kQr5czyOXdqaUCbvbdaskMf7wJgYlkchcK9Hs
iEZE7OQvJNjLkSnXBw4i3B870/qbCbqzrr9jfdOp4n6TiNab/muLlgzMYMR7nCOiV8pAs5FcF2tW
jv6a6Ykh2LkQumHqQn2VFLvFG3Yl02Tg3ZOymoMAPAH4gLfBBBgqaSOqg9ckOfh1SY9CxqxDXHN8
NGCN2+pra2canl8X8sVkjVDwkTewk70+tUz/zlWahCD5LRPXByvV9UmeN/da1/XfgpLGLzWhk3lV
9Z78NtJ2nObIvT2OOF6mqX8n5AeyJNJTmeBUE40K32fwJfRK7xlZy6cZEgHvJqWaZ+yFz3MEgTn0
JCp28G4Y8ch/kAVWv3/4UEIY9Cx+NAVuEzPgEqJWbNB0wKI/se3s/NV1YhCnz0QzCw2ltF7opi21
g/nNinv4Nm/0OyBEGC+UjY/168tlc73usjhX12/jf5X+ESo785KVwa3ObfoQ2dmshYF3QQQks+7p
QwssN230bOrR1kGw+6tb8T0SJQK8KtRrBelm782zVUs4e0xRQObTy9BDjdujWi7rDKohc2popTDk
/6UOxYUszeT4W9iK9UJvUXyWNbYRplhzlrKXsrlyOqU8CK9FlOoSZNgjBe5p7dkaAY+ruz4dfiAr
0ZR3bOLuwhqKCt0Kv5tXHoIufafvd8OZDKanWcbFDp69cbRdUIDCVQX8UjtanrxjVeoEhBbOidhf
3O5WmqJgiUiEKK2fWZzCejEBsvYxnbrbQObZlMmrCM6zS2c0qXtW+jjEVzHjjWJvq3rx2as6ZbDo
I4FCkSAun2419dkS1ABG5Dc+BRbdDQ7Q3o913j+rfsk1/CdNJHAM+FGR8/mYknzZ1njfsm4/OUhe
6wEqjWFRgZ24+roTI4Jt7eM6r79puiBNbj2JPJrUfxwdoI+bnAuReoN1RXGkIPsHaZM8lL+dH9mS
ATzym41+Fq002364PdDnIDw1wcprDGp9i9nITdCCMaSf4oSJQvfpFLiuOrEwMak74lSHkpUghnvC
dI8Ckv8eAMer1sX0bBokmG8TRW0AxGJ69TS/IG8XZQS+Ny1lddeYOpLxDVRWwWn49TR/R6UkTMOt
p5I5ZVLhEBb9Y+3ekpxzVtDmP11DctoFnydESaTgI0Fp6P/h4PDL4BLHxCzSexZWo3ScyUROQhAx
RxPdWQne6OVTUgaZSGHoFztsriHRhnBN3r1oY5inVQNBISygAht6rM5z9YYvNjIPwGRH9mw9Gbtm
Ej/V6EHyIrHsg97HAirUCF1yY5b6632Q9mfGQYM3yesa4eA+5fIuL3etpP76+JrgF3lD3ts7AE9x
EGB/pXPsD1KsAHVTGUY3d7dCFL3MkeNmHClvuiQ1M8t4BaTh9fL0WNKkwmnym+/9Z/dAChDjTwBr
zn4YlrHMGSYzraRU3t2rq0rhdiTMpfmV4ypxXsfXZNw9vFfKzvpwUgba4A9Fs7kYo+XHxY6b6SwA
pNlnTjCBojnUVG0Zk7sf5G0hqlf7YNw5EjlSqLWPaSJfdL/ZGBfPujP8UMb0N1OFUtUc+dhdsrdY
xpVX8/CJQSS32X3GQx5/sESq0RcpYpaFaKkFGqK5iGG/OEvuBjV7/sI+zpdBXT1re7dTrKae22BG
qVseq8p47wT24l2/j6XQabmbEgpECRnLy2wM9UOS5Ut0CKGRWDZvE6pSpQGFyd4kIk/YxUavj8mm
wNa8mupQZ0eYu24PbnzYuQzNEN77yS+QCRh40eJ/VDzes7MKJhehNY/ms2lSj6lQmYUI9bBdVg/s
hzhOAoQjELE2mKaYH/6NTh+pElErzmIC44aX6B82wPCKPk/fIvsT5P84CzZFqnwVdd6GTJmY68ZV
v9ZtC2lAtOR3P/ZZUZ2ibLllKvn6OUn+qsUBYvkzg8+HU6bwZRlkHbx/1BiZBArT1ohnTHG44EA9
QAIh1lwFzx7ZAlH+6+9ZYTM+f5sImKGHdp90ltD9EYfu0CCWBhvmRxpOq40SID2CmPS7m0QrXlwz
81P/puhNEth8UThGYebE8M9kgELnSs8tATivO+prOWIbXUcRNXUkzj/NaKS2otgct/0+YBp0pezU
vnaB3AXuouwWfQrIbjTsa8mWQnqx8TIhNWkM7xCGmD5R46ZT/TOo4EaIaK5p5h8wYzag1JgI8S19
Sp+WYJnlXrIGmppk8blmKhRVC6BRSFjUAOF2/oL64Z0w1OFlykPD16O0IGRpgp54BCHf5a5kwWKo
EGIffRUP0hfPzoyWYnMZY5zkIsTjF952r3/iq/WGtjNJ5RT9R5wIJPmiV2ZA4vN1QUApNg+n+X64
kIXgy1pjWZoFMLEC+vflqkbXz14UJ/Hk9Pr4yE0zmobFfRGgi7sCpOFMBkBDg3pdVmtgrEEa+NZ9
BwqJtFuAdvsyE6RtFwVDcWC37o5SrJofFfL0mhixJ7fySdsaySz4P0eMhl0Iuzg43Ns/WnJu37ST
EWRvuN1+xewHd0D6i9Lpk20yB4lDSspPahvFe2BtE2i1pJEcSNNtpu8PNR2fHVGU5zQ0FSlCUQvL
ppwiaLhQWlQOonSU7EZqdCB3cdQd1X7iBhbBEp/Hm0kocra77c3LRu2MZK2rjdOsE59kZ7RTGEb1
WA27DHrQhn0Q0/oBHsON4egVOvYm5seBwPvHkoFTp4zb+5rNOaGzHehQJbdLcbjjmeVoFWaJQljp
4J5o++oRQPe4yV++YpMF7b5mXUjwPX7TGmI+16pLVpcBxnZelkYpiuLLxTRY3pJ/jiE8nS9WWIVL
PG+tYfNfULM2s7OULXLi685XdWJZBsSfw+gVsr6qIa2B8n9l3jjLFON1GZo3LR0E5pLzs9nt4pW0
TTSJKsdmweQZ6jUQCPl0iGpLg1718kj1a4RQb2g/XNadlZPJj9G/d6eSZyttuq4lbWdTyqnvW3YR
Pg+lUExwbW+3nwX29vCRGFyLFrIlWIuO81dkJzh6ig35hMR9Zs/zw+l8QoViy+EwhE93Q82ng/68
gAt8eovlwZyZIUSs2ts5rTREKppfq7kZrpYI63WyvATo1Uo09uoSM1TkE0vgBORnjYuKuV1RZNRl
Lw+efh92tzWQjWd7wFD31NEbbWSU6M4cvNipN3Kn0N5AgCnGqPCZsMNZamAHA5y45QdjXhoq55Kx
sTj2a+GxaP2xdvWXT5CamDhCzB+9sgX2lbf5a1A3RL/yP/Fz3CPwQwAJDzZjBNeVsZDj7WlnE61Q
qQdYMcsQdInXzPpoH/nQad+vYMUp9IIlVEQm3IVx5yxD6aLZRRfy1gXLqmVXH2ubYUuW83ApEE/e
sh72u+qY8I7AHE8BV7+ld8lWL32/qSOFxXrn878A8ZmAXRsIiN4em2rL65t89jbR9SRbEF3Vhdq0
gCqLw0vUNBylqJ/CZofYdYR0d70ZsroR8vVMfSjJMFjixenroPOIyJ/6/i9+uc2Ut5c0iCBsNmvk
EULEWad8iDjKV5/kh/pgbSXcE5o5gHRg9GvG/P6xC1cKEji2VqhpDuibo0XttBsqaf+KdyaNHMV1
elEBNg/eDGi1QeiPSlO/U6LcgtIKI519NIChBMQiIkFLMdLbPnEWTuoqnhN6yFyS1T3CmKm2uvZ5
afdG/uQ+Idx5SlDQh7YpUcuoz3rx9eqdTwh7cn3LdA/2dhQS+h88YVuY9WoJC8azTeQt8uUQbeN2
4SELarJmUf5bSV5pRbyZ1BL5+2jxkqbMASg6kGBQ9uiuTJz9x7YgsK4rQMf11mDxKwvQFS8uHk7F
dVn1ozn6bjflaGSqIuzEv3XOFCCqbZ05MtrUjUocR3w1wOx//V2RGZ16SPBcj/IUV7zcme3NsZvw
DW5rRpiISCDVVQXJ8TjOnopHa3Guh1FH00E96lc7KkYQUKlwUMczrlkG66xI4Xk5LfgycJUbfBYq
Rv+13OhpmYyS0rUAbPM1moGA16FcYhKwUnV5yKFmBpQlx3ZW6lujw6JnueKcCuPhjghmA5rO5Pmm
HQGA3SCEllIo/q+FRrrBOwxgdL4FoxX/m0Mlei7MVDWDarQNQDoTagQ8xqEaxJwfUERSEOVfOBrq
OdpzZuGXmqcygQP5J/exzdTCMVcysyhjDarjJGFRncAdA8I2mg49+7st17ukoPl59Smir82ECwd7
xGChwvjjL0qlDO3juofbafLH/RNCEHDTmOGd9eRHA5U8f2G1bSxIK2bQyoed0oVj96Si1uUD9C5v
UkOFg4zu9G72YHwXfuRrbNIGyZV6AnX+J1jQkw+s3RS/aKUgD82VsQVNExV6oPLd1xEVoa42nogA
Wg25TbMJS0CtYH8Hg6Tt2Q9qSODjbMtC6mQMFaqWycAS26J76+wqPswEJI2rCukfUOxGFyLrTipG
UtSYzKg1wH8IJw7Si3b9sAy7TTlWSvGAFwfhc+5SmlkwNimp1338ReXIDOsvuydewrnff4Y1/Jg2
7ZgHsQR1KWA94QT/r4hmZJ1vIo23KQe1UZx90HMA1Bv1mnack9a7NIu7ap9Wa8StQtjt7++k/Y/n
+I6BPwOzaYd4tv0ShNboY7F4awvKofyQb5wlDvlTTWhQO9jsMSr714B0Y/3i6wsSf/2sTXjZtIh2
yvlV0LbcGjFMI/B6R6/7jnkmK/p8rubvqI6JpmcotElVg29uk34cuSbi7pFpY7cG+O14zlCLfr2H
9MbulRr9cUi9/C7B3yamXB2iftZu+8g4oL1gCBmcUV09yHGbJwCTuGoKVneXTra/FA7WBu+bOfMw
fEt4tBlQH6lONIL6HxD2s7m7RwTwKeyTCfYkECoAURJ9GiWpvOey5pXlEc9qlhi3VpGZ9Ym3hYOD
QvfAAkL+zSI/yI3avpWJ2kAe4HA8kz/GjqBJ9YWHL8IbeJfr1bpk7YaJKpcJ1+dIxgDH9z/2kCc9
DeHGQaMCFgIWT8JrSroGNVOMUtNZk1+kei0ZBvcoO9ilC/3jsy+opNzuOWrew5G9S3b8Wt3G7BHq
dvnq6ntvs8l+Fe6QDGziPTP+1GD8Whqpw4uI/bAotNkAS5vCwTktvBz56iilbrB1iW04292BYAAT
jVSXpuoZ+KYwOYUwmXpny8fRGhlwbzGpLEh27oUX4+zrweESVEnPnspZjnBPYL7rq3/sI6sVRMOe
w4E8RpFsY9tTp3bE7RFAoIqsaP7Nu6F5ocj+mAvdxo9vULBaAUTSSRow3U6lMfV3TqvX5crfNP5a
hXQ689vrs5vKgCaleeZGrYE0IATPWBS91KL5BANoLL4wbQWvXH3A8kySC9wuLO7Vkh37Qba4iN3e
Wvx12c9jSi7tSbz4NCLxe09gm+gX7rNjMRWTs/gBsSPkJx6t6H0xKTpgCIejrYNfAfjhwZqslDQo
X1SXLzXmGwfvwO0gL28FGy7oVm46Kyx7ZvGFo5MPN/P9D0kovlxMC56nuTHAZOWrZINd5pWuc7Kb
QSx70JXpwS0vRpyONidZegGyWjszF2KbMvaJgFAWe/4G13l8R1inMFas+Umv4Ph4CR2aKW1cjgsz
Eq0m/KAM5SNlz6i/bxei1oyg8ipYwbXLoaLvX7EOLY8MwhlmNN5uVusErfedSEnBmTPVgwdTpf8V
O2Z10EuClz9Ry1cTYjAhbxHYrhbpmvKaipWVMOduud3pW0ygSld2QdNTjcSh+GQdOnEy9KxHbFpj
NNpfwoJOQ91LeZCmnD2Z53fYKmF2EbjTla1yBDpNVvo4j+MViaxHlSEbGE8syVInjiJdUZOZE4TL
RfeHlMshYgBHZPUbXuuROdONMHyCx7bAsSyVronCgV70aAKR5BOgzdLG77CtqV9xbs+lgIzZeG+x
nFX8++Mqk6dvatfAs/aoYd5rctnAJHvj8SFYtoDxE8BNv+3G0OD/nRSDrg2XKQg2vZsWKPlz/2iQ
n7t5/nBMhyEPSetIcIdNXyEtSNCtO/XhyjwQoYyO61NcbK9Qp5EzNs3F/Hha8vTSPRlY1RESpecR
1NvxTik7/pU++Zf6gVNbIx/CFK4CreGPilHCWs7L21SxW81HkG/WdsCwXLeaH4MkPPyjkTtICH+G
0zVpsJi2IhTooJWgpWeGlDnavgMuY5QGdUX0ls6A03z5JQ3RWuaG8IcrxrVI+Q1fzHt/Lfd4k4EA
wflNPyQrkUhM0p3EfHIHsD1TeImzOvsJfO7U5C7/ZwgR9UKCe+JahtbcTcPFiKlMsOxND+e0F9Ff
maqTuMkvcd01B4m9TAHiXDNH6BFBAwgCqnTID7uxkBq9FzP1JDX79GTyYTuqPqBEk2bckk7Tmtuk
l1p6Gbcsw6RKbPUWcY46ZHwVCcqw+ay5gZoZod392eoZkIx82XjmHy+zWUQ0TfuKFdgNS+vWE74R
YxiX+UDPF4N3ZStQpx5ssZInp+EULlwr7C1Y3W5cVCU7v+HdkKuo189/6MaIq6/+57qxrtCdru49
BfsA7FzqoWy82aqF3LFF60611PhCXfW/irMMWZTH1olBuOJu34qLEzcG5wIQ5kRnBfikK1Og6cu1
Nov3KiRXO2cn/PBkjDjRsOFRsfWoa8ecY+GxBiVG2KILv4ny6u2E4DCtlRDQ8XyISuxciR1bGKCZ
P4AC+Pal7Rl0R82HruGTWK/c8n62el5Y92y6RLXWlImwhVgq6nKbRPrweqHcI1WEQZEVRw2up1Ek
F43Sutib1xr5/wsLKm6SNXC4vdvfQtPqPMHBz+6cQcBLBccmlKsUEPlAyd+NbqzvQvsBmGIOYxY1
t+dkYvdYaTWnBIk/1T/ztix8q82FOgCqdigCP756Mpb9xuotnCnDXO+SvE+PRU2urT9WMoCC9L3i
L08ao1tiKkno/173RKp1Jr+9/EJwtiupDIm4LVZzHihpOe3QnxRaknk4K9tJa9vGQo38slDK1+Cr
xGgRCC63HOZgAaSFavv4cSUkMjiTUh5XYXszd4NRZeZLc6SfqNmKoR+ocYaiZHRr5feI+hX+UKGA
+FEPYU8pcFxbv8pmKNi0OUKI8ZYSu/+P0PP9igjib4weIVzm6H9hHM2hcAFLWe6IfqBjBBIX/SaK
YblSWWSLPyjtGUun3Az4FVAlbOQlVvQcb88TVmAU6+HGtzYyc0t8QlkxwhEFggHYhgqG1ddW1zYp
tHJZtmuAaWxumalVYh8mFxxGILHtBPiD90UxeWTK+Tjosh/YtnuiYAzidn2DzXOh1pRPGPCApcAf
8oSwkMdaY0L5/uhVww4tuKSWY+Y6iQU9E07B7MJwpp4h8koXXmnv6BBcIhFiELRewH8WZczYSdv1
sBLJtNWuwdLWaNdZy5yTWKRhvSP4X0KZB+iKBnZ5gWkBie+LoXyXC0d+KU274NW4uszQM/Qxa3rx
QeXRq3MMdz9xHIf3kWD4nBN1gBtjM6M0GGect6OpBrp6XatwjBP5j3mbh5yNqZ3pZvVMTYVDi3XZ
mDOvD+RNq0dMjHvWVuaGlIa7ZZ54XAM34vGmXy2T5eSiRdMXzWLCcSCWdgxlAikZmBvSMwwWOgpl
T8q1V6aq4QCLZFlVk40AxmeGdpQD2IAs+kYVvW8YmLmOpuT76vCAJitaJx5+FVMOBeOS29+EfJnN
CTZENfB9jddB1P4LKKuDgFUgxBh782HowEY0dRbIgeW6y9XhZGeXIsEKOPOM1Zqxo6ih/IJueEUh
666mmSAAY2Krr0+whPlnxHAo2WgdLy+CwurPzZ/ShcVm/pVBWkMxPAMLvQuyvu4ipEfOBTqJQL0V
HnF8M1XYEr5IOhyTaciec2fSUi1iusUOlL9JL4k9BuZv9IH7mpRCD+1qkKK6SFBlSXn8cBqMiAtu
6mFkXs66rwM3sYlbOqS70c4nr8fDEYhCPyDZMNdZZWYZyubLe3xRZRPzyyCoOsvQKIdArJVftmHx
Ku1zi17E46ocRG0pbiaKkIuKKiAttQ/IWHZRX36da9chKMfjXlQy6uKqDWg4FWktX+0dGSqT2oKH
sh/DgDqcAY6a9SUfHUIHOsWnILHzIbS2s07b1yi5oYGhQIzirBMUOv7xUE18wQJOKq8WUkU9buDx
uqwJgeSz7X9p+tGTMviWVOQoyy/JaEbDnqVHi53V+vVwwENGTk1rzzZ84dvPnRoqIHZiJEJd0QHa
ns9fSHJPfnNn9vOtg+e8NB70Wdkdl1uHhvM1cLfoHO/CPCMotI4LFuf53sk2Hy98zp1JQYOU2FkA
+/jjX8M10/KHvRyyjBIYSUoMdMCSmJCovNgeEgjmSu5who9Q427YUBKZHMWkff6CI6JJkf3D2DwX
GyokaeN+zgXPhCDOyB24gvDDlQQIrPDNWWpMr3+ElWso72rYr3NJr/HtTESOexmvgx69Xd3JR85H
HM3Pc4jWmOyguZkZHA0HmF1W/VNlpZo/y/QC1fDThvAAr804FuRh8ZrH8kxC1DabsTbNURurZXTY
oDWaQ9WtOlW50rgn0n+eyKXamLn9YiV9vZEsvrffYXkvzExiVzeVH9+6ec/Yhr/3mNq+ccpn4reZ
vMjT44n2O3gkvqTK5sixuBGYkm7xqhTKbU+xeVkskY+Bkh94pRbzy6oXtjwOsi/nwVQl/543XLk7
QBivXVdx3yupCAANrfAlEVzQbhCKG1u0hGo5HudjDXIfZND90X/7kcdl2jfwgFTKiUnrtjq0QFBs
QGZoCiJAdB2KYrlR0NdyEIGIOlQOzn6MMxLN0npIPes6oGTL+joBEkwTOdsIbX100bVtpBQJzKSS
qO8BTf3C7UkY2zN7Q32SenyApiM77mpzNNKRS9bM46Au5S9D9SFJxXYwJBM2b2ynpbXYev8i40kF
hT7PGi/D4aUnaw4xVZSAqKOdxQPZx65sxKOkeeRbVYtq8zS8MyyCGgoAkSChFC4Cp3gFZimU8CWq
QZhh7RZcQDTgDOTFa3QKPlcTIXtNAm1GO0T6VAAVzAQ/Dt++mYXJVVbdjVHRYAyxMH8DHWhibXqc
qKiMrh9Hw9zS2Dc79eRwcu6PsnXVst/KqUxRmOXENvek6xylQvsZeb2GduR9wPOWJPwOj9Z/0WJR
taHkFUFCWUD36iRoWy6uAZg4/qP+RKhJvC6N95tiCPiqazf5ccucgi7EnZ5CN+7uw6ic9UzGS+jQ
X3KpFlHUhL36yLTmAWUxJEtU8sP+tIwrBs5T0SmaMSzI2eUrUlgBDRanGbZv9w8balEWSGAT4OTt
SMuBcr29hMZGjtzefr1MHnkgJea9wNqVdLrZymjs5bW9kFcHhkQ5PEMm4WUKq8cbwcGyNnN8DbrH
nv3M96AOvm1QO+dJuU7uXBcFmYefIYhAtb4Zm08vzObDTq0ZkpIwyOYW1khjwM5X+KfAbSLAtHMh
C9SaOiAVX7IJ4un6UC8kxiZ64dgjtfw+mCIP+6se3UuVGP/qflNlaD8lcG8juVfJP5Nu/WPkJ9H4
rmgeRfMPX6xS+dXZjuN7eXHhOwuko5/6gl3HSh/MUOP8CcaGbfz653jFXWJ6XkaijEVra5S6Ocsu
I/kNHU8c+wj3OYOuwd2TB4Uc2/ErXAChUZY2ND0lFFqHxY2uUbWQctdTaQ3jTneAmofHsoBXppyx
FCffIHo9rsOYRgdrJ9LnECkk6mDuUYfAwPeTWpZBxIN84kMDLlPChvMEIEMCS9JVYlaSzz+JJW7d
eNmGc3HAK8T+S6q2GdWUD7e5yuLCugwl4K8mPG3hDRFT6t9iAiT1JJ1GgzONgAcfh+y5Fn27tt3h
0nP1o6xegQWBf2WoPtvB3t4z6QLp5GRu82u1sAaGs5mKi3AA+PUocQygF0jzRlAiNmYbtT//hnrJ
2PXFdhxM17B4ErBmLlea/Uj0C4J1MRzridKwP3kJXAUyD5h6+D1q0i9L+KgOIyTUa6mhyt0zLpKv
6UbZQv48rGugSrDEIqpXtE/TRG0cArkWFAmoLh7xPDlWnwrauaO67m1deOCPzuiJOjyH2IzVEWB+
t1SOApxWSoV6VX/gqkNZOdkAwAIvJYCJBi3cr8xf/c4nJGSzNlI+6Uo/s1mHldTeR4WQVQ8jvqjp
h7V9gvrIDUpYXhu1fpkZt8CrwDhpWC4IIqUgz4/qh/QndzD4HnzIb2PM2Wl0UGCZAE4ZTzdZNP0l
RSOxNpQc/onrhUR7fG2+VcSzzysthcik72ozFF04jyKMPPo06Ta/uHITCLzTUH4F4KLR82FxnzXJ
GWczPaxWUqq/KGg3kHjXXjoy77Q5N+hCEtHXvn/9RNujVGvXf0U31GK25zlNrmx5xDfS2E3W0JHT
AkKST+5gKlpYlVsDfAxBkDmj4ockzIKrNOp7hOPb57XgwDDDRVrGSQI33ndfBQHXyP52vYGrEK5x
hGcBq1M+dIoj3CeEOqmQg1Z/3RDi6TBg2NHLFVM3+TpWZ9ALcE3b9/va9P3xsXyhNCiyt6gdrGHu
TSdsOLRE1Mha1p2z/2dnVzX8s2U43mOegEuS00M6Rz/RWCwJUaOc/IPd44VR3aOLkvHeHirofOru
eEsUf34zbBERSmwhBotqmNVrEdnE5mJjnMEndTsr8SrGYe853m23hiDZ79mky1LGHjN/HSJGboCN
Qq/zkR9Y2S/h10IDaszFcliWW+IdmiHZKeF3RusgBDYJYD+J3NeW8ztZOB8nrzBOA//+IMZlmP16
6+2QU5Me8QGM+nWR8Q79CVaeY9v0ZCoEBCWOpUACGR+aTC4tINUMPGKEUeBpNCTg7UIePBMADlJX
yrecxZUJNcR+kChkxvF/rEYlVXg+O8baW3YMpv+CQ02Oq9Np6EMm4HUBuTWMiaDVjVv95evWOKxE
iybadhgcN144bTCzjQNU4BGYn7dhbWP3JboXpejZKeg0P8rSDbROni1cYJnuL1t+4wcBS9USWuWn
RbSWwz/xoGSyireRrMDoJEZB2FUMuToPOKscusk7uL0aFaWjmy/rBQz2o2WjjcYETJMFiTzRIGND
zY8gO5ydaFiHVus18Q25o82laV9XJV2aTih/p5ceYVJC0FMH+k3MiFwjZ6AXVuSfITTby5cgIZ9d
RSPDvGO07fZd3JwRl/lnM7QfC/8kZtG5GsyZ5dbyPuSOkmGRKcS7UzHlukXTA0n/leSsStR2adw9
w8Xb+7bW3BfzRobwmCk6NcViRGy72xw4l251Ub7RCt0HRy0XB+3LuTrU4i5NbFbZOD9k1EEAu2h6
Xth3P3zwldDPy5hbE7esD/9POuSNFNSPdqd565w79SpUBKel3tFDQObXa24udmBaqn0ka+GVqT2O
MHECX6vd0NMMMjTv1HKY/Da3l/UbJRHdFUo4QJ1mvzSL24wW6RyTB7xwimcZSJS2XWJ6dIncHJ+1
wXRkSQYIVTXXktVfsqPlTKh2+SXAk5hx4NrdwAuyWcUgujWXzLAPr+15dknMMXbN10Q5ZC4Fk/t9
cWJuz0EyvWvis18bREQc+phbxceqEm30zzcPy7uea5nOmD0cFllugmIcKJ2J8sTrTsSKA65LOL7f
+0uZX2J/4ZSwuU/ztU83tjr+LrLcHHfwAZwYx1UidEhCCKaS6CUQjT6X2y1jSU6I6rtg+8bQa2nb
ANx091ZozrF7xHbqZr7Njlzury5m6SIQVZ1hw1qqsqUQcLQAsNkpzdqc/ZjT3fO0b3KdlxhVkTMT
C19SSeYCdex9/tvztjYFDjMmSm01zNiafyCjkpq2/ECAdpBpctuIS4D0flHJ93L0+Xymp/SlvQq2
lnPtfSVDkx5kOfQWx89Fugv6GGWeBggWVdGuPprVwS1X3x8Dd1wNvQDy0Id1MiH8AuV1+SJ8VMt+
BKt3+/G7npnUzHU5i/ABEgg2IAkAVJYQQGuZTItRzewTZrs5QclUrGr7HgAjRPXlNT5m/1lAu2s4
0Ef2R3aImi2wuWSPOSh1H2blaVQjZGFo7ar8pU0ZrXzS6/+i/qfJ+yW5XywUxvBJHueXTLGVZW4H
Tw6ag+cRRtijEBM60c9ZUhFLoyZzk1c18np8XuournkeMenljZDYah+eupXMGgIt2RiyMfdwtFxd
0+TMToM1FU/0PLWWfimi6uFzonYMygpchxGGkiT21Bl7OB2tFTpMdOPVIq5BnjcjyKlDCcc50FBt
wVvZTIX9R295Lmulaq+mMo1Z46H1MOIEehQYCfYOMf05wE7wr27RZuIvuiWF4GPwWzQ8z9xXz0Q3
pjmENtUYjeSaR/VOcoazKLCI22PeRDK92tqMDLhcmFipgZsjbjEesnl6JV5yMQur+Q87grOt20Mg
XI3walVeF3tHQ3BGHDQyn22ElAf/mOAvW/kmge3t41QJ7ff4+wuJ+soEUSl47DcxjcoaPALmswAV
3M2kpEs4yRPM+dwVsQfHKKMN5abL8Cbo8I1jGM2TXw/JwnKykSsP5w8R+cY33XHtX5ye2+jQ76eR
BjTeu0fS4uvfNx2oCgAmsd81a3I7U4IhYf5dSSkAtAONQH4EYukiNhrFOwWlp7W5IDnrXCZPD9OW
oY5MYsBHsculZjDj+axFTl0xEMQAS2vSvOQJEZdbdqaOttUjIisImAZdg+tqDv93PW1QQArayOTW
wNYSJZUF0c+tpkCgleMP7T7oMflTZOINQdF+cl0NbQqAVrSiucKSGwt+LsWce5fqbjuLJMXu/V72
rfirr9GbzpPzceHorTY0cGBGHVELapz8rl0Dwp7mJhqzDiN1O76iGIbP6vjNX/c1CfqkosDUlRKx
V73MXrvyTktJPmV+8pE3vpATUqa9qHDE1VzoGkeYV9+0awUFcdpWoaa4CYzEMXzUzQkqrfESE9mQ
ozI956OhsMzN15/CAH8BZVK7GKk9TyyTmsYcYFPzLONjA8GjNqMCMTd2m3IheSuFTaDZZ5gCsx6J
raHbA2qgr16colfRRez5q6ERYIPByReeCnIHD1FBHhGkTNavMwMMw6GWKBNKGkr+AB25PQTLzFuy
gNZe95auVW9sVuxWs52L2JsrpcuH3hU2Ul3wgmogdvt1tt8OHA+l+Lbmoq5fY1bfAAMixXNf3IF8
vWDdbgfJ0WXqPpPn4hd+ptPMDjVTwJJw+dn14kaVf3tjnd43lyxmHNnA3FNDOIm4RT2vWpaJKFdc
RDVflxE4kEAcc6jJ39GOfzKAYsiUDPcQr8B1CwyeOzMdmZkdgPv8hydaZhF9/XXM6FynDaoXRKoI
i9XT3U2BXLSnzdrvQYgKODUySTCXSE+bqul5+d2Z20/5RR7w8iIg0DjF/Wwi00YhnlszZmj0ebIK
kJJJIl27zXKDGF4vLXLaL6snpp9Q0SgCnLcOHFiI1HYvO/6dQRvigFPGWl9DSysuqOiaYhLIA1Gw
Diw0ONhelal5/FDUPhn/M02SN8yOd1csWCBNN4OlEBBW3oPZTnz0h/QCyehoilT9js48DhawsX6G
mbrpmN9FSyJs8rhZP9su3KnwC2w+upjInkN7TiC7aWvXPUlim2cjk7Y2Yxsys+xwCVwPGIYdeD4g
gq4S9Iv7W3YlNuEccSyipy7vxp4AknW3yAJsTIIzrF2LDzf231sazDPLgO8KerGQhkAGWXgcIZMo
boQzSEa/pWM84sxQcoqEC1iQ6OMOBIEt/Q9n+gceqgWlRaX8uxslMn50Ac24bSoEg1DMcTDHNkJ/
rxm9gxJJmw8c4G5nd19b3UN8hVfgy/j5F8qVr4cwyDB7PE/BsiQGvzkOh5k/wyePeJwBndEY/+9a
eBwIvy8kq3nHgvn7mTsM6KX2i4BUVG+RKayrxs1nGNqLrdkA1wBUhQibo02LMzlFZCSku5V73NcN
xhO7KYlKIMWgJ8JB7bYCHFJeUnA6PqSYrQH3IgSRPyHXl4icF2bGZxM18ftCWKCuH6kcNeNt0dcK
7v0HipShE+IgKGa0ESumumosn9aCe3CqTwTVhJhOxnoTz++JpmwrMjo+dBrpzeHUODB55Q5xjJEX
EN4f+L7//vPdcb3KsDeftFpYJJ0n/LGGN6seHPiFQmIqXIDL/nl48MpG8N5cxwsDaXhrDNc5GioQ
1wDxKQHnXhrXQsjO7o3Tgn0qwPztjBIVpM5hayJaWwm0uQtv1sbBs5dLmuihmAV0q/FIM7m3MwRM
nPj511+/Bqk4IjpWyaTfckaL/1XT8bSmYpAz5UesaMHuftwstkNFl/1HQELUHPcsFD+27KAjkMjS
UMQFj2IVAvAo6ypyzchgGNXViOZ+TNMFXeurmx2mxV7OAyMz55Fnell8G0D0ICPZublcSaS5/z+q
QWfmlrl2bBEunFlvcQ4P37wP33a9Mq91wcjpcFLhkqTsFICcxa09aZzwaUk6y/uHTCtAa+Yq+MC4
ZgTdkaTxsqKWCCb3o5LEGQ3Q6HD7FETn471z98o/ARcS6tEVJ7WsrsFou4zjsEXaPy/PEVQPJZNu
LdwvUJFI0aX+BGOr50VubUm5Q3Pg0iz1UuMAPRasmogtzs2sZKZSOXTzYDkNrwdaob6ThEVyVV8S
4p474aRa5U1CvrhxxvmJIteTA6RI26xgc1A19Jn/Sx3K5OBS11HrOMnonim4FVe+ng4VNCoktVRL
DB9cPoaQIRT2w2TX4Gz3pARcNFz3XWl3bUJauIR1OvDFU58gKQeDXTKLrnFodixeSJyr8lvtohmp
GfnhH4bTsqY3GxHEz8N+rUO5CNoAQqskUepc8fBECnznlGaHtoZXDFhpLDF3vv5WkS+2+IIn6PM+
Wakrjws64fpliL0ZeAunlbI16bR/VTKFS14FSFEmhOExXK9uiodPl9wclRrPVKmfM6qGN+TGBmqU
IOinZI7J7OIUd5o4Zs3fQXkS15upOUNC14IdOnJXW+ji6hxKQgRNpE4Fve06smLbrPh/USQ4+Ies
qA9MyshARiQg7zRdLg60WlliX3phJRIS0WSCgIrl2gh61iB79Oq2y4rsg8wy1L3BZqTCHcL81hCs
Ehu3BI9l+hpWQAfQvIcOVaOqB/OwsIMXzF+QhmjkpMGocmwHh8ti7J/ZXZJJQPviHIrsZu8twS7C
rd9W71vuzDAUrvOFPAJN5VIg6NixTTbXmVytAWvyeCTyeUNfzzSOqVdNmp+ppgmdI9VVdPS3e+QP
WNx6PXXJ5tkv77b+9I5LiWEMYN3IR8HlV+9JQmbgaf4HpO48foFlGY8gAkgTV4PaybS21foyZ/Jx
LuLvsRs0O6L9EoU9XRFVukKvQ8WZIEBfZhfnElwgXnO9UIaGBGDt/FxgITAX4qwKespPmsoAjOJf
NFXsLztgr8/8a7Ydsv2zZJo4TDx3cuzA8YZlmQ+GamPwK4ehY4xX4dECZ3yLMaL7zK5ohW1yhVIE
iVPznLAPpGaJR+4eUoerEuQIICNuPSwTBW+l0M+ZEN+6zGx5EnSpZzZSmvE1h33isPg7P7Qk0I9S
t8R2kpVcEgUB34H8z7iu98PqAEgGJi25NFGPGmEPf7hm69Sfyh2INXxW7r3y5/wkxAc7w65crfOE
vn3Tktk2/mQ+9IANfBiMxTqMohuzdFOOJIElIty4I2RC0LZZ2uDsw3fANyVC0VLJFtXxnA7liTTn
PTJAqBAWMG0ggmnp9fQBXxunXkykUGt3PxBJceef2I19PCCRPbfdtiWdsSAOUT8FGr69Mvp+VamG
ZoFl/sAplf5pr9KKI+06t9oT5KXB/lK8orjNYrmhoFJXMWlLucezVenhn/HhwSK0T8rsATtQRBo4
JS25rsr1VkCdD4aTwglgm8jcfnfOn6ssyX1jkmc/gfO77HMk21EPyJBlW9e6mg7FzwImFW/yXkEG
vUKzHTnYzpaCx5wbmxO8IGrvNSJ0QX4ko+k4evnXuAOxwDdxjOk1HaNZFCX3DRtvU2V9mqyxZHLx
Gg6XAqlb0r/8mtrYZ7IWMwVylwtyiJmXzILC+0rKSKk9y2irHt1Uw7TeOgFmyiVcrRZRCqslvTzV
GveQSo/wZvrU7ViDJHglHTtnFrfyLy+ZqzPS20jf1XfKPty0CFWu92/2TSKpKGqrQ9A2rr+d1+Vm
Ut575La4rAGOSE0eh1A6u0PzAtDJxt1ct6W+mMZIel/1aHCU3oGeXgXlCO3F1VOGrQj4nj5a7hfv
iO9Sg7Cnm8R1FAUUVf0Gwrkn3VK3FWD1JWbwXo+t1EAJfFlv7Eia/aM5To97wxkWfDu+qa3CuQpj
ZKyK2cWhrW7Co3KuWk9wpIpoA+LjpPj8ANqBsFZFQVvgnKXcoidUk0Jlozgvu5K8ENkiR3vndM2g
9picN7MvHcIY8F4ZV3Y18F+Tkc2XfvyVlIVgHwDLsu9E/pAeVDsR/4LHOl/epPWLDtTyaix5MwoL
pDZxrqrVUCKjUr2kniCdaQa/DmQ84jTyLoUN34y0PAe4BkKa2He2zGc9SSSThkL4vdv3qFoK046s
jWilKhK9/KlBm0/xeJYi9M7paVNMsHbwy6w6l9H4p4SyWVVue/vyIJdFyGHJg0AOgSwu60JJou3j
AUZDUoRIsGIijl+JCzFLE/vutJIr330GP3Dwt6buGDL/C5riSdN3P9Wl1/hJsxF3+12U1GdpZWcU
wdMzUB2RtJ6AIeWseckk6phIO9dGUBoKyGd6nGjwwF+pEk2+xiX8JxKGQd5Ws8qwF8EET5YUNqxo
uOnZCB22u8gFa+QnT9ZXxJ6P/C7TndBI7YSNPoR1iK1s2g8jZXgw4j7gDVY/L2UzdvbzbfRsoq0M
4Knh+k1S464qLE5EKrPq6vpzLkO62S9Mskq6rDaSrs6U0bOREzRH71kzpG2VS3plJqHw9eteopT7
L8NQJJSbZ8pZ7vxMh0+0Y0rdslbYXdLn0t3uvKbWLqkgJ25DXcM77aFGhW3QKUfzNAzByyITDw0S
Ock/TwnlO4LAMW6zr0kmUH9ZLzT4q8/O6Pr8OmWrI/LSYgyDFfMAivolsDQK2uryKjojKkCr5TrN
BiNHyO5iElUIN4/Ow9wHhH47ZaZjNr4h1A+Che36Mbwc5qB9IKJbUSKZN6YsYoW5EiPyqz7A8x1w
coYrT4bF5kGkYGYW/buBAOUHkU7iPdejjyoKJ0rGb77rofjWlhpLVxS8SjxGjaS8qcnGOvV/Ie7S
cjis3u7gNjQvKWVlNN94mxexI4Sc+GbfL82q2ke0teAoHcqBDnu7OXbH3HiBgjeJxLV3HmiL4iOA
iR0aNm3rANVRd5A/zD6tzb6NB9kA5O0etqAIrqlho9hIyKqDxgmoPK+YDARPss1USFJb2jon4K08
eN5j+YgXumaOS2BfV+q/1k+en6Dtu4A395ur2lTHTxm3hNdRENr6SNAsXmhrh/Vzpiq6trNDjWtY
/5fYmdM9X7K2hPk7bBbuJonfybQtGDBy1HU0iuNhJGVycPrNexcinOW1lPyJLhaBj/Uu5kMkTFCJ
fsvJAxKPJqNG5/GtPW/rk6kzr5VmR3GfCvFBUwjWcuAEth4Fasqz4ic9/Muw83t3DmrZqpVylmTj
d1QOryMPXNpGCKU8bDqv+OnvpegQDxqLLe6mu6O37rcsdTPl2epI5Cq18rGCrtGezvr+TjS4onZX
FHSUvv+08JOzrw8RxMS2UfEYxfrcbZWEyiBc9czPcUESpK2iT/3sk8cQ6hzs2oAHn7UWQSw4HSPR
iR9WdJDW62M9bDPS8T0oA7c2TZo2/n+A4G1reqsfN7NIp6CrD1s8H2w+MXiKVPIoZnnBMcZKPtu5
fheVVtbboSANxvqWN38iCRrI3sRayS0ns0LuvsAO28V50i4J2zhI5dyY/gVZwJpFNQdz0yhE3q7r
390S6vaE1cCU1FlsfeUFiWXXKNDmJGim9od1S+zZSmnUO7ilm7mM3UxtdXbi2QzPgLJOyHpDsWJ2
IgB/RMcCLqBMTeC3HRV9X/RU+vZ7iCCRydvT3xsOIb+0YDNDiRWQgqA55WsepvSHvTX33rPL5mMk
c5sXk+cpzfxR5DvNzyK3uKz6D6767/epucIJz57n+Jj1Zxc8kv23CJxR8/dzanhtc5f/dCachTfc
xE1empnH92mwQz3J1zA18CXMz2AI9zgskocNyi+wR+xVO+/Wpl2CgWWI4i4YBO8HtsTKWwGMqdvb
CyJwOmb/Ebap/zfpJbqojsDk74fJSZDr1ntMNUW/jWCUkjsvnxcM1sDDwd7pqeKfrlN27aclONN/
6T5qe6eEmMdGNn5EF+XiDydhpIOiwlrnYnm68hPXul5GQOC46FKZlUpAXAt8+8pRQwlCkYBp3w6+
zKQS6ve7coO8Bg+NIH1O5FxHL0QJcJ4Q37QM4NnT6kdQXcA1ez/b2nw0qsl4ezXoCajU1j/KlbZ2
V38Y5VygLMMG12cVEYUxQ2dwvgryLHAQZzrr7h9uiNnWw3sOvZpJoiheFHyjEGaZ714O36EJQ/fJ
yrEWQUO3NzLe6FXsDrGI1643NWm3cC7QDhQ+c7YKgXLF4ubaUrJPCGNZyZwkpfx3Ff1jLmuCVgXT
E9K5lg5SoF2/tUNC60tYqbd2dJvo6W1SIS6GXHXHg+sChpp757rhyRbf52ecX2pCAkbQxbJWgvf+
AAvhhcyDUv/jepwXUOTWgn3iwRDB6wfomUEKl/7VfiO5XIUaJGUbArMe7PQSpsBBTtPjnGLAQPUP
YXgYCwO/KwOdMbdagn7bCjn86GxNWngpR00NJMgPl9iGhXImipwo10ru64K5ifRLXUSuEgUD/xED
aMjcIBS23VrwW9Av+Y2DExIKjxlfHImfbF4/AU+1Rs+nDIY2ucRwJOYhStir943o8IxdaPVC4Hc7
aueCCZA0uZ3kpNTCmPcsZjAmJjlr1LLAbUj5Yi/xs52cIsbuBee57p6OOsrwSvDnxZgltfX1mXph
yj7rzkcq0meahwujeu557fOs7sVO8B/bUVDcHrEyVv2UOMfk9JurUL64Jbx1isx4+PVT8vhzIv+k
x0qOdVXt7K53fbgabh50LeQP4pQbkWy99F8MDbs5duLLAeKywDDLSkKLANE02JhayjdTmxy17cQp
hGTQtGEaBE4qaqpW9vmv2Kpr4FFCwNhU6/8FUczCMcD4URNmLlUwN24es2Dp0n7eZNgyiFL5jbGt
yGKVqxgRYkQQ85VoLLXKTZjv16VjJhpVkJ4A+wTZ0V0xFkJ9jjZWi6lQl2BHJK1mC+lCvVWw+gN6
581wt2hSurbcA4VIbiViWB9I8sznkQsX5VOcd3oqkasP/tPeaqZlwHa0M5Ce31T42olTQxPPxcE2
kAddiyhlCzoOcmKX706KJ/Z/7OBDL+RoYTa0NdcFGFhcc5+RGgE2IUVQY1ZhYwHf6Nz6Dp1a8IeX
FI/gF9gLF9WVsxZmkNbsZtsghUeV1Ixw5reUE0wlzMfIY4hgCk4ZUzqLZ/6Rw5+VtK+1MP0S/puj
YbnbY/FYX14qq+iFEVv/h/wDdPhzx+KDVnr2K+yI8+Fj8i2wIjEoatzYKGc11K0laiYiEmGM8LSq
4wLIQP5vXvbB0GdIJkQ+Ul+ZJAUyAOjsEb7ofxOeRiNRhz6oKm7tcW9skxKZ8S5xhqe/jpeJr9/C
a9BVzimTZcjV/Fsaw1L4UqfYBaSSVKVLW8SasR5wPJo6XJTqdzZCokZ+hrxoEos6Ilq4vXxa8hSv
x8LDDSfjar1vVEmUnZRRalaYo7kWykZiiclXcsL1UkU1pr+a9dp/bDrUeuqZLm63k0GskxdvmRWP
DhN90BoffE+ypG3KWLG+qXeDwkjodYo8b4X8db/7/wd5z30k5ezqaKm8C3SlDtCIchAEDUjDtyiy
WqFq1F4OoEzl+8oxf1EHNEH0nNQILnR4AvwUDJ8WHcrAZ4JeXZY8eNXzZHCnmq1LqKaDJe4PzrUY
lDZ2Hx+cN9r4pqd83YMEuPTfzxdv13K0F30hYgrnNKdIJDxHrnGkKgE5ws81haxYclDwHEwIrY2T
II76LGYx6fX7wCRDIvZGaNZET2n8zsKULIvJEXbgk4POo3n/Dqjbd/HJGgD7z4CVjtrrhmFZoihZ
UDi4SH8K7LrPHqNPRWxAzdfh/T+KVM6BDSJjwqtHelTaZ9KwZibEiKP+9LQZA1zXa0qT59ye2s8t
0Yop3NdzNjDfNpkQA4/KLAqZXy+K41neHPmM8CklCzSlfhAtDW1q5tH6bQ9TZXNKwha+F3pPxot7
49YVi/9vJcjqrp9vuoN0RO7oizdaEDJ/IU/CtwRYyU5M14GoG0xi+4HJKvu7MBtvZtLWuNlfNDNQ
0LV2AgQz59jz+vnq56PwJd+XmonOtBrx3Mhm7VEuqW0nBE1iRDaBEfSO2Kyv72bTOwwmBmJ3agpL
ZDw8Z7peVzT4aLspsRaqo5UVuvkMTj8vBUUtbkE1oDcIDDH8NVRp4Pecrp/rOG9UiBRCCqQhul13
1jXTxQxmFgaNQEd/CxLc+PcPFswj0lT4VGa3VU7KXpUDcPUfIKySy4Fo65/jJYQPeQ63eueKJx2U
/0grAT2gMH9HZGRt7ZcNFbosst7ybIrdVeNtjrkT0FQS52OFeSpETm2LDzMXmL81jDOycgCYorVq
jFMmFmIshkM/EucUifsx/OB4RWPSUvRIeYq12ioIf91cZY2KIa3toBNoxOOSbiqcMbojWo7LMMmq
WgPDv/Soa3cN7g2aArn0BgA5GtrGbgCYHl30gPFcwoKHlyuUYWq6YFBbHLUR4tDjXezCFevS+QCM
pfNY1m7r66MejXatHsm5eLYJIJl7dWwhFBNAKdt8EUIv7SPjGueEpXMritro8X5Ys4qXj12pSm5u
+HVPzhpxn9M2nNs5SdIN1i00c8xFS/q8IAyNBKrdl8AtyZgxGPOWiSltHcqVtX6by4VgtgcegNx3
rY7RS4CBLi+G2MgbCuumKkUbpZMPgfPn8WWNjKXj4KPk8yplOYEL2nZT2nFMwZUD+kxqwPZsR/q2
GUUoXMIZbqWd2tjSjhviuMg1DwxL/Lupeach28e9LjGcCcdQBJYOw8MwPdjP85E98j4rXuRuX/ug
wxFBm1P4KCe3WtDXqQqFGj8TtJFB/FUirE9s9MQbkIXlE18rqmTxz5GLt0PGq9nGEznkJeAuzHrj
HSaiSpbmlKa3HmEkcfrHAuffrICzcxvzYBib3Hx0JRRc/8g0bMB9EZCqJZ0g20dOFA8gnGP7AU5L
m9L72L0C0W1g+aWMlIQ8ZFjhfm77q3Bm/YCa0vYSvYYgT3armH1qq52ry1cU0OU7PwdWsfUg6TWz
/a+Q5WfhUwr3dSZob+ihi12OJpTn/geTwd5TB9KQdXdtvWDtbkmsJVP6Keie/BKD/8CZv5OipiJw
DTT25rnLvHVo/5bfwIPeLyce9fkDWBLvvw5XPm4ue8TFp8AMilv8Yr4SRqZUbYxHvINxGc0wjNYI
IujnQGnDpw1ke17d+LuluubaBRSKAkN+srEnYj88ZFNBOFBHgSB036Tyf4dE+4t02tNjb611HdYC
KwRPhgXVDMaoZPSc9QWiTeIPImG2t04nil9GJMVV57wGS/AzMBkoELprnstcDypyGewayTDAZas7
fmwfr1Vxex5u7oV+Wo3/R3E/iIZfLazQhPmSB3rUR9Rb0Uw9Blg5D7cgXo8ll79YHn7b8XtL2oAt
7hbqAwqHYv2PB6sgMDjRVenjf29S3ZhbsnET2zf9R51z8mpt6c68HAOEOWPb8DJnXz1U4rE1cTmU
JmgpDP7RgLdY1fCpMFZwJmrKbFVz5cu4fGHPVmbiJb3rxTy84GiDAGtck1uMY2Hh5VOeDrYqKYvc
BlaTmiDbbhdigEyzv6mPKmBdBwKD9Yx7vmi80oC5MFtUwxa+bEz/NpjmDpK1tHHwptFX+B2Ux/xf
42tcZg09gFPfhhy1AzwOIxMhHoA8hKvb2gqLaMUobMeNdQbGu8AgBbWRdGCOnJu3VJ1SuyXLJh5b
zVlHfH8w9HB9SN9jIFA4jGZz3nDg7kz3ouQlLji+75lMP3YZ5uRauRVGYvP6XmObD+4HpWC8QztT
wrVg27cizrWvcLVylIK8PLpwzCvr+VQVuSLwOY2i+FtJfJj1hXQsg9P2dfZqPPSfcZBG3yoESoFV
O2fKYaDBdxLkOauZ3/iubToDzWPZtDC7VwZG6fTt/rx/4b80uJq3L3HX6d2SStUjZsFRcpbGQBal
93PaYWcY4/J75bIbqSy40cjTH2Zhc3hB97HNFm0BlpQytUoP6gT+mgf/SvnkE4qyFVfagpsVzvYD
YIjetoJ/HD4bEL0ZUN+jn9mF0GGG2lzhKj8V5hZAj7/kEyRiUEaPIvLSENFTDwfGUOyzO0h2RJbn
8Hx0prrEaDA46+EiSzbGYG6sJIDOG4oWx9IB73tc75pcYSyymle8TBJdv67P2k21ABG9Jrxckm8f
taOqfJHYyvH3RvTyIdx0AOMaAflPXj4AS28duJZlMK947La2FE2C9yWfR2cxHvZ0n4pq/hp8gr6E
gDEKFnVPr0x+b+k65k1ERhzaWAkyn+nhgFe8AQd6dw5YjW4rCGjmAaoX35WtotmQpSGaV+dg+2RS
xzZ/WUiEx8SG8FXaJSWHenM2LxsRzJ2amgCfHP5omPC9XDOIEvVo15Ai1nEhkFp45C2XTffDDOfc
6mMXbYFGvU1h5CNRpmXEwlrRbXY19E3RJvaVr4YJCnRPcXQakDHkjggSalEe4FZM5pa0+R1VEYab
ZaEfd9snYjCgFFWZ2ZUZR7cedT/tkUSuizsmsi2OKBQnnwxFPKa7hNVe7LzDv6p/Fs/a0cPFy/ks
xHpm4xtIi4fvv16gABhu+cBLmfT9g1uNiWxqYjVjhFtK4XU3qh5ksB74f5zCReU5PtmBLAwEuNko
1gOjP3qXrM/ogyVlDgeuqLiYOABwmZIeslRd05/9dz0OXTVdebTsloRNR6aM4QpxAUEGdNHC7v4r
F90uKp19rtN9s/Zaz8PPmVeApxtgJMeHwBWalkk2FVWJ2XkwQN3U1tsymgeeT9kBvWz+kFFAM3IO
UUXNVZRx04vCGTpuI5R1hHDRqGSRGnkIPrelJMK//Kc6UJBudf2ysCr8TzGntCUwh1AIVMlaDxUt
ISSZYKKgzpJH8F1TalzQ/NmXZNRYQzq1diu88IJvf6C9nOn72QPBDXsDUoOcrjSRp8kCVnaGaHyG
cWed6XqjzpW5/VjciBFkh0Jd8MrstuQC5yPa+1kPVx3zh//AALxj39bKj7wvHI9tNyeWhY20tSIO
upmsazfUo+8uJItDr98U15DCMJbLjq0sfrm9o+TIGGSPdGzweE99TLoXlxun3DK8gP+kPPx7dwxJ
3ZKDCKUG8NqljcgqqITgk1KbaBw6CoBS5RmMu/3H2w/xdxgHwJ9UpTkh3/c5nM4cM3B28JMy23J6
w6J6jYEg03rl9RJ8gtNE9lZl5yNgtVdvj0YfUduTX/X6HpyO1vmgqbEZAPriKlk/ejD3Los0VwW6
znwANmY8qZdOHP7JnE/+TbjySaDVC4f4YNWdtojg2svaPACZMiqJExY014gp4pXbfIZcLQueI6mf
k0iDvxd1Q3qMBJTuO+bj01r/OkWNmSZOCfSD7y9FRpLp0OPo6TSFqAjTMKHTQ8nZsma19rAlUXAE
zfJbED2eC4EyM6+4DQNSmVEO1IEsR8fMMI9oVbm6QjW8apSFEVMOc2H105245UJcfk1r+GI8Z83O
pfX016RvZ7zuZ9XLSZU3k40aBU/NqSvsZKQmjCaOlz7O1/qIaolyucnKw8UbU57H0qJn0H4RV9YG
G43R1Kf22FbrLg6hGVJI5G0EC5X5k4wnI/C95+oVQI0nlbqcP/mGxBlJZIx8AYUVEGMdrMJfRaMm
xELluFVwG/8blrqx9vc60qrrM7g6t3Com+KuwZEgj+oO1xTwEUQdAK8v2uzRZ5gfdosO+VnWqF3e
uEURPZTb4Mp8zzRtTBR+wYCwemXiJd8SDoDIgnJ2+YAUJa5jUuvBo6W03h5mBqaVL5Zawp8YvyTv
qdXms9Nurd4uVe0MbmFx7eNUIK6BKGxgfnYFMpQz/iAKT9oY8ZXnFvfd3XySanJ4SrGJ2irnGbMJ
s3HBpMKAAblMuM/bJhgRgQn2YO6XVHJYT40YnqzI6uT/8fC6C8PtlBND1wBI8YtbZmDlmqpHh9IN
tyX4kMuLeg3xZVpRWBzHV57NrBm0lJ6V4JrHuDmRWNgjwfZt51eudOZsg9Ap61FwE1jqp2Y3n5Lx
M5j0Lk/5FP738/c087kIY4shO52JnAYYiiRF5+rM4S1ltjaTZj2iNWVsdXPNHF0AOXEyxNJkOkKJ
uAMa5z+jMm6hVADwAR91O3fcTD/XndngKSkWtbGkM8ccb5+RUKMwwpA8z2PPm7QcVoB1KtJ9kK3h
xEiSpGO/+BjT70/65/B7s9/wgBfE2Vk9RS8mQQS5bqC0E9o4Mw6NPtuYWRfFV4jpw+VpedQ+Jpla
+Q655jLHURf2g8rcJ3rHcL05jbYXJOW7VJ8dXQDWspMuHnZJ4OO3KwS1XQ2Ro6qnXTvOHB+grhP0
fpBpYFG0bbySzAiA44v2do2dISXmiChu2aN+R2nauVIutPQqL29b3wYg7+kUbF1B8e/jIXzPzdB+
9BRsJ6J+jiE7KPwn+2ej8H+HyVgYqQJwabCqOvTc5Y7otO14ADCNH/LKvVYWQwxL0QDpccWldSYG
ITGrYVpK0lbsD7EY6FYZucNp/no+K30SWvpi2AhbXozFwZlv+P+HxFPDHWNUzH2hMiTBRuqI7pok
X8nuuOfTjPj7kZn66P2hw505lheIxOBmxPVW1JcyBVaBtTIK9DwepPP404xpHFhJXCqTZP6HKs/0
x+WOCHv86naP3chdx58msv4ISjV/+DOE9K7ceGzPPesMw3Mmb2sMx4F2HNPTIIDfq7eznNEjbU6o
qDq/1UhmxA4ZfQkp/ti4Yls2sszqU/MT1CwHXnZ9FiHKidAoD7s6I6kD55Sd0WuC9vRFKt8LmXpM
I6hJ2cOVM+DtYLNwd3spg9FNuyi/Sr273+sD028bh54e02Nz7N+vSy9nSAcxSVVwMTITgqP2J6bT
Mmg9AnUpRt6RkzcI84Ft4u3aGVaAzIXQPCzNfBDE5lSlbZtLF5lUT5/SPb5gFt7VuHink8VvYPUH
Fm6/I8BIEWV/XWUgJUm1FNdlWfyHL8cAlCxekux7pHDfycLApMU3dNqPfM3Li9YkuAaUy8+gPVpZ
sjWKzpYUiHH2SkePQI6/BLzBt7wTgBELjLKJqZeeguxAj8Yn7xerj1Yf+I4QncfVPRoHZzdvWeZg
mzPVEwq4aZLebvk4lsRYrWEC+Fn3e1QnloNS2pW7wISWge0uAkriUh3ABgKOEYoqJ3C7Mant3NqW
N2EvMtNtrxzBNb9ZV0hP5U+0SfTIaAn5jJsqxyAWey89E4NPEQup1MmGuMgk8Q7hJHYKSY2p4kgv
RZ/RtaLDiDV2rbRRrJYeP+eMyybhTxIDSpw0vSpXiFObt2N9rzCycAS2RDD1tLb5rXT91Qf+nNHG
NhKjGKviqXNxGojTaWWJ2U7fV2bH1fIhA8112IwCHSE9u/mxKPObwn0OAYVOaYtrlEsiu8UfS041
FoYqVF5hJ3tIfp3elzFwqvoSGVAqxI+Y/+aole12lp2ZE4RZ3ioMo9HBRo7VXnSvXShXb2THP9md
hQW2gt4+A/khoKJHnOVMQK1Igz5kHBapA1lDEN5HBR1i0AlAPfmKz9V6qbNTc062tbtDhX3yG4vh
QaNaF+dTxGVf8lq/zck88Jm/iO27PR3gpoZBZxDP3mmxFefDaR+d3jRoaTiadDbf7cJEWrI6xY7L
LyYa/gePtFdfSezv8d5oeVzBImLVnb0AJnRYsmmNh2p6XmemD7mVNVwA+hNN6lBC6/8glWuNOKmP
JRg6BkYU5gJnks8ZQaTdIJbK4E6Bcc1w7EWA7slI5iEuj61+IjvvOcHZbo+ZTvy/8QpV1lp5r9DV
hB/artAzZufpGK+EI2YpFW2s77oGynf+b9dRJ7Snz/jb23GtuzyaeAQlI//ShFn3dTPbFO1PW8M7
tOAGime/tWDI4TXS5zZooadIM96BTCGGbDWWxLjBbTmrgGTJNfKOSq4e92p0rrkxl8yuwFmm1Xs6
APqeL/K1ULkT4cxS3//zJ5zulKg7xgzEhCc1QlL19czg+FkwgM3icsDywx6xHtW/1wVvj7Mgs+/8
214FDrDuff7dwFKeIeZop1Q7/Q7cuYw/eBCFzeMACMR141TVUeD9SE2GNk8aInoVQIa86MKJLIWe
0TMBGIQm4sFNWwZ97G8zaNbhcVP5+qKz7JI7OZeYHZXx7kerecVhsZOJ4isuzlnrvs1uxyz7fgLr
lSXbWRa0f30NACrMz7q0zdexnNucbD/ql8VQ6MFR1kkIHhgLkkLZljt0wfnMgqGfpznbosgAIaii
L495bARAqGdtFg3v0I3I/4Uw1IEmD3rO3ZmbvYgReo3jurOmor9qJXQzRpONVz0lLHeYCyGLY35M
cl37ZGo2v245OIfiIgVKb6XATbUScHCeMnObXai1DoDX/dze0JmvGdGjUVbHXy9HZDsA0hGxx6q6
pKTGo8MSn1774n2jh/OX7GUsTGvVun0HM/8Anodln+2swA91FLYAq0bx9ZTTOFZO9k9dlbBnxXin
mK80m2V25Z8apRG3Y5p99AHbsk1GRZMIjcvW/CCW2ZfDhiMqRsbF+Q4Sblq762bzpp9ATryEcLrN
o91iXjXaKyHm09+EXWKgg4JsAqYbTswAdr6KEzkikz8Wsarx8boAHC5kQ2/BybJNiiF2dDevfCMI
NnS78jw30r5/GK/KXsusTCZqrXeEFv/KpNI2ixmfYjeusTmEI8nW14PcayD+G7pGOd/1mnB1XaTx
L4fD6P5QteyUbZz3HtUvuvrk4Q0CRII8Hho0211CSqVfnIGKSlNYYlDgw2Hm06RvDYL16su1GIIb
2F201CxpxU1tGYtzHD81ADXO5kOUQ/9fJP7mqBCAdcOcW/LVEbZTC7kzyXJz95pRUGNlLJ/QfklO
X+talyh7wpc/naWoHh2R3rlO40JFrwqnmWEKu+thvhIyKxR/mEW4JnQapagDMnq17Fxr43eHLoNS
gbphuxwH172tfjJ97QpKr00sYdpyYpNX+DXwy6NJDBA3YdmSZx3Ct4SU8xGRCQrjenB6yAxkx92H
T3ECzMNISDuzdyFKf5iqcmiiceVrpDvQZ9Ku9jo/FBYgYceEHXYYPOyhOX8QXeMfb5ku02afH/cM
JWlTMeiY6lvsX4vxG0Vlvf7+SZ957BIXJUnRoOuKq/TywKk6M3voGCNuHqTPe0WZtcqmlYBua0e9
lOCDyXgQgMOz45ekSITDZNke3zgoSqtetLTNPho5R4P77gJm0QPk0MU/CHabxwjQc5516ElVncUi
8cN3r3LIlY0/UO7VsMchWzOpd60TOQaPwstZiamJUvtdcCM7BTqwdz4CPWr5TQA5Kt10tRKf0Us/
GJnnUT2HT6oT4Ud+/piZ+jumIVwaMaYG79z8v8jsXebpUB2s3nYfpDRBZPE6el0SE4Y1CcY+6mNO
zbhHjMgB7y8hVsVfN4aRw0Nob1KF8afuZ0qcde3dEhw1MTe5oHtoAJoVutmPHuHjZ9V3tfMqb/D3
Zm9RkWiM7wnHaGP2pPPnaQfVsAOgXaCu+ZTDSRk0vYJrKv3a7U0pF+8oHFJ0hSjQWrIqG8nCG6Ld
VYPq7knEAOCYEkKxPNT4Ir5MkNN98J4ePgm4KUK6oKMZEQVDtzN3o9UgGEqbbEYDgy7/yZIvUJHX
7GnZVGkPGPqYXaGcytMvFGENKrfgASctgvVwRIRCv5f1xkOTMgT1nBSDQKSz24Dlr51QHeMOha+r
1EDJ25Ga+xLn1bpMGaUmBiJQmCHeVJ5bfi2kOhj/G+gC3w7B9u+6yKX/NqzCx2dmLmfwqvHdcVZM
IVDvegJzJ0n4mncNAE01SoFGZoH+Y8noWjO/cW3mL2gfE6ul6+QcJZ/ZIkcJBQ2fseYifY2HcRzQ
X0hrIzocbAwzXHENfvN3OGEXhGA92Oaty6HxIcqZEjaApYKf+yyaKAz1QMfghjm/dfwmakEGxyqA
yKiNEj9w+ihuw7kfdPDICwQSKTUXpiDNA9Jj2QBPU09EB386AGgQgLnZobM/WSE+7UyOiaUSv1fN
HBgb2E/SIBzTzWetepAD+tCNv9mPR7i3qXzojUAHai4qvbCSh60lzVjuWbNzn69KG6/vt7EAOCyX
Ggx1C5D2+U9/f4ChI9cwstKloe9H9qH7TlyJPOLzixwEOWEQ3c8qMMBtAXJ41aflurvJ/Ux92Bbf
ZCVbCpA3yb2G5MHY8XlmlHIhrehTokR0/ul8BmB30tZnGko+9QMo5+T332KGXIX9Nd/6nMBU5Uzn
2oYWXUNw0mVKiLD+t47wy/z7pAJnL11YdRJcaLtVmyR4Abv2ajlhnx4kmZzl3xTYkeaYnHzGDCYT
LISLcERmrT0MOTcz+wAgiXsmepr6d0y0RMzlUHs/1PBEjA+4EvmtNvPZ03ASOhcUoWquZ4Z2TVGM
2PWVi0F5eIEjswvdUFvX+HZY3hU/skfy4wtT+VKcxeXLExuGKwbpQfM440GUYTw2jzdBj+WmPPRr
FpLLIfNVZvSxj8mkfPwCuU2lDZXKa69fu0bdoJOgHhIhmzfZNR3ZIG1OpLcT6IzVC9IfCTXT935X
ScZGWIesa8BkmzrhydHXiTAWF+Hlh2FpWKqmESR7TYY7cEaOp5V6TVQzWFGFfnbw110z4XkJj5mN
CZOW2SJ4INlMYvhuRuasTrJgUfMPsX8LlRRu6MNnyxT3ZNWEeMcMVY9TvNK+pDHRVO7KDACkZVR0
zY/nkmeVslvc4I/hyANpe9kN7vImkkncs0iMyhzdkB2+kR1F+zA6k+id+tWUjPl8IdtR0KGK/wHX
KqPBUCR7amtfI/mPtuFVQtxrHiYuMi/PVZhdjONg0y41Al6dOTehnqGhm5QgwyNFjYBg0cyWEmlO
fOEGj9u2f++Ipw0ykOpQ+vNPT+zysX2Z3KbdqDKWuUmyqZpqQ585qqcPJ5sCf23bwYLfhAY1v1/N
e7QTo7sYQtcrMymm3mBbmMVWYE9+fZYZyez/H2zuqcT0rM8Gt93q89pY01vhnKNJ43OdAO0zt5mc
gg0N5Nt+bCMPZ6GkMkVs8yWY1KR1KW0mhobXpSZyohCcu2Ol4luSMfezVDAsvTBTBRyk5fjjfWbA
6Jpy3/yjvDP5C/7EN1Ir4p6zeUs34d+xu/AMmDIqOd6xjtBrqHSh7nbKtjnRsJbM4eUQF0I3HaSR
KI2/OIE72ZCophCSlotDF/OZACrhXLj924m4S0AhFw515m357dpgWhSHLeX9XL8A7q+sTBEdXY1d
P6QKN/6tzmggC7PzsRLw6ED6CavqUnhOWHNpIq++f/eWcJXhYTKGkO/lul6VPfe37UWuBx3SVV3s
2RZgwLRk0Zmyyi2DSh4mjmfekYRwgyXZxtsejxD5dIppUwRASPOmmgmIgd27zYjkwwaZ3Ve0urrs
cLWpzAtOTuUMZLfsA3PPvb33Wa/ty+q2K0XvTH+uF+2qoiEzeppRPNgcNmb9P1DOglwqskUaqzpn
67BzsqcXE3MiKD8cQuGTY774xsLAJmkWrjZMYNuyu3+IDEl2b1ePPVsHYmVgNs5CYoOLyVnizpin
aLsdtSwaEILoWFa+Psc9VsrhKJhOTaJviMPKwnWB/kPO7PEnuda4MZjKqprMPFWMMCNd9eH5lSOU
oyGmrYCvzQgw4udxkLDw05rJeWqsgaxuRfCfFSLrQCedI4GT35RvS+ijgoS2F35RsPUcAeWLeAeI
6oa0b25cFIHtNWUwDPROl7GofziSZenl67if/scxotqJ9RW/w71B5lDd9Nvtufgx6nKeYYUBSovP
wbPyZnU14GezQf+xkoaHsina4k8133IE6ueXXf/a3VEP14Jf2v8ZcbOsRNIOEyl5MWpb+pph9vew
HjnA0U6gH/p70kO0PPpdP3HRG39YIDOoWZeD9M4B0WG3lHlr+7R/hcGIhrYcSOXbvB9vxiIcyvim
dLNXJr4cvYI5tKRQiTv1ogk5OenLSkn+09vCt0PvuK2EZCv5i7Q13jKfLL1ixNE3v1QgP1Og2tbH
oAiRJ0DUhiI/3GHWlOdb6Qd5eEOLEc9X8wUI7KvIwN/3U9eRIMr73PQlPqZVHw7xM8xKYeNImc7L
jN3RkA9suxfpWPi4njhd7ozrqzR5++A3vIdIXmwhbChoV+vdNL9KLxZSfjhHEPeYHcoS78Yy5SXh
lRc/yuJP5MfbR3xjVmDALOX1acDJnfSDC18KRmYrEnbvWhkjc4B8TF0BXngtvI42iN/vf/vDf74E
GzDkPO1GEB8nEGTfiDq4ayUPG9dbk52d8XzIojOOsc2PUpEqkpJAnHFw6Ljh78xn3FZHdxxkQQfu
0AZMOu61IvB6rz9KdmFco7DdGwmiFOZ8cmmoXkJNtzWmGnYTTq/8ocku1qlOTcDdQflJOtBmoYEO
p/vclPeiuD36V8hJ52UUzcT6avXt7H8pEcEZkn9eq/XYVclLZVUicVWQwq4HtW9QQw2/tf7wlRWd
p3erUsH+Lu3mXd4ilbeAUs7XlCtwIsGeFyeVkq6grDyvjJdH1H8YBUT3YBskbt72IEhJdjyX0l+I
+X0uRk9mYF00VJ0VXq8iS6Y6knHy7Tj6le6MuGtaWlw4ymeujkqsBDbSu5XDVw0KEU0VcvtJk1hU
SDsdhT1cdGY6rz52NEgjx4xEMQkOT3TCHv7/+uaEQDEkifa4C5wWIVpdki6fl8x9y/37hlQo6lkD
UNQ2t0PKMXouO+EBVesZ34u+iJjtW1fmcEsM5Cs5C2lJtkiLKEAgDP94VvX/fa87YeScNEyS/Z04
xLYOSGALiAlshajTKNwEXtedWhYbIWvKoheMzX93nQ2k70f31CBQ2e6wHUw6CdJ+TrWYH4VV6DjA
mMZVAQodssCWOuc+DTu4Y30nwqgtBnQrnMNq2JIfQ6an2cGJfY6kwpBytFJHcVtcio65hzsaWW20
23IOpUiPOTRWNyXBJsX6Y0cj3xZkhgE/IfOxy0yxCkGBOlwUEJoPxw0xt6MJ22GD2r+UDo3xWAJ0
3+cpoOMMs1BifhOr+PyfmkImf/H/O0bjw3lz+kOTG8qu78DuhUaqeKWjA5XO7EPhuq8xfH7RENvp
I9Va8Z7w7Fo0TDvKfdyJeGbjzl7N/TyYCM/sWW/A8HiZg6cBJvDctW+TJ9+6yvvCA2UsQyCgLFwz
cHGZcMZLc2ioa5Mc2xh2XBqIzP548aZE7vkG6GKc2nqeyl2tX15Yif7H5wfaHdPUamnT5tglrC1k
RMut07gef3uENnpUsEmftHlEhmN8AmeX6JgjhHMd7cfF8apH5SxbPP53N2QJpqXjaF9ZJUelov76
Mzu1kmivWy5q4u8AP7fhuvcs98GrlLG3wVW0zIZPvhJj2R/DYKDScT/oSa68Of0vDTgTRpVUIr2R
cmlcTzk7d9WzFr0G+hdqw396GGP77V2eD1zJJvOco0hiAskoqEqFWWweUxgb1JaDxsMpEvx/wP0p
KWSLd+AGGgf6uhIppadSMjpANpZK4Af0cYOFONr08i1aKp5tPbEyKgydTVgW1UQCKLAak40PwR+X
9nox/QUrV6hgalv+CdcMhb+1ttKP12Afb9E/GR/xDlXEgG1GWPyI2uU7dOzxZ3yErqXyqai23xrl
iHrLsOcyc8lfTHGj27i73ZMYtBmKF/ibmF99bL/rPzRl+LaU3297BcyE/ldLWI6jzSw9Ai5lE8Ut
o7q5XIW2ZL+ZfluYXxBFxU0p0otHEZIBo+4b60Q8tq8beKR3/mVtKAjagTuPNiu5i0CXnwC1VX9z
61lNuZwhrgQvFkDoP3XX27hmVBfhBgfXJrav3AAASvokrcTcawOlbFR+97BFYqva5CQk7qlGmsPG
VlEQ04Wb0GpMTSyuXm1XCp28s5eRd7V4sKa//q3S2KZmgFWYcWiPL2VBkhrYV/k83e7p2zcVPfeM
tNwrhTxOubaWJDTFm0WMegVSkK8ZdaFXDAxciMr3zfmKZHIIpV+aeY/+uiNBO81h2xS0QOts51mf
TjYNPLH8lAy5TI8rEwPCb/ifXNk8svwhHwj15vrz9G5XY53MQ7qw3LvjEncoDKypJbVsye5Fbqdr
+0ALM8Er+6DdBSqVAIxlK94AW/Q+17aLnfrCf+qyBsWoGt82iPJXa90eHZFUEbffANszouip0S5V
svViGazAHdiz4y5HAOEVnaXsebcd1edbHSQP/jE+Ffbo+MIMpSqGyypYxF1JygHPub7DQaWa4NSg
tPr6FGN3F7c0J2PIPs7oWe0tCQ1az6wx9e/NVjguiHvAAlal6HFmH6YDcXFftQQikQvO58fhz5sF
taPdmns5+38/NPDF1w5U5Usw8VGZL0PV8vCOrnJr5FxYz8uqDSdN/JAZ5upTV6GdCrczMHKOwgzm
lE7sPJn6KIVN49HlkLDQJ1rtWjm8Iqpd6mH4+OJLVGvvRbcz6q8GYBi/ZQVuj242zZgsJhg/apsY
KEMZJNgxTtBulYDv/z5VNLr3dp3k0KHLOky1aJQKKEhop31Uw48a5dHpTT6+nUZ3Twp01XP/Ca54
UNVhwA2QkSs6cBokfRuaFVoVcuXdb6sdEBxx8Zv0FVuSrGMp9pug6NxsquRCls7LCY1teC67eQYz
Nv29RBtGR+tb560g99Gr3k9YtqY/7di69Jvyj3TmyTtn0sBU88wTfMqscDeZgo6zPKwWSepgBUWn
QCEYHkVYo6D5vw5du6qn0oZdUZG8WxFtFF67Z9mQOuPZA8UzYaXJ8BrWJL5GCfdybJqodN/5oRhg
Tr32ZYzD1nm+q4bY4NURW8DFYOZsw8wgRagF+j4toQEDhLgFWoVnCczsJTdR6sM0mgPgOzx6OyiA
TygN8pIW+Cd+WSN+Xs2x4ed37CNnExJYnPJy1WvQF7XUSFbKdTrPgMfQMduoqEkkkXpVBXt4iqLg
TBcQapXoWiC8SrjhrlS1BAjdcxRDHOc7MJzblrwE2Wq9MYOILPos0bZohFxNJelNrBZKYnmXq0CY
0XQ7PyIWIV1qaPfHa5kpzOVh1SCHQb4zK6gDeamxORLQvlqWLowDPHlXOylpIb6B3WHiymAQjkgp
vBmwVBJKJDgVHHDuof1+5wmXvVfktsiJ6GuhWGlto86/aMiwTltJpYjIWYvtkV14u+2XsQ2ID6NL
Ikd9NsPaKX9oCuYH5lEWRBCOvZasb2GNo4nzcmS5mz8EJZ30AkKwxhWelRXwUo4CIKImuXvvO9o/
yKtQthgklAW8Zf0EKMyg89pNez1/h7RJ6wbQ30PwyDu8a17sraHdg0R0yuf5nS1XTiYF0IddHnwO
JJF/VANedook39Q1EGizhKH8oHST4NMOVzxHB2/W9fSTuF12sf/wh3r791Ue/CAWJC13UjgMj3E2
ESprPfr23v2odGgT9J8yySKLvCy4HBZsxPoqHrOvdXEJUOQKdcV1iXfzNG4di5pc9TOr/2nm0356
ycV0ySeW7KwZ9XDEQKEiYOxhMEnubkKXRT1d8BhELnuTet/X0bn+XNtk4+5P/rIGEt52t/Ynpvc2
JwmblwnV3fhcX3BaOd7g00xL0I9aixqLNhi2fD4Xd4jFvBOcgVOVk/NcgWHOut58pi87rudrY0rl
KQPIshf7S3YFoMKQkICGPAdqOcqPRixoIDlpAs4xxc2kKCgIbXpXHw1+YMHFwA5rEVf+IQymNBPh
ID9F8jvPspMQjoKkp0alBz254JAjLQ5BIlLTZhcB27rcd3ipXZ/iC3BZGJ4ia1Hje0qdjaFwm6HB
5x5kbc5ZAlcql6NICFq7lYH+C3PcMAzr2QYMpuanBSXN5U0cKzxMEixkvLexoMBBkZl6bnzvz7cT
ZOkgbjL4PS+oJP2zSKa2+CQMq1df3L6FrIhvKIR4ge5dMqme22oWE3F12AoCvhOd5iwgVKs2grtU
IC46XsI47qoCKW5q2xulihNAQiuFn9KbtsKYvHriTtNXYqwVzyEwpd5JBdb38RhsT9tFblCkSTJA
TQDxHe4caNXuVsQusBOkM65yprbfKaL2Gx60yxyC3AE3w7qLLV/67wAP2wdnE2JNjv/g69bMx8Hn
iTojyQxOSqBLcpfBrGodwtN3bYZDKimD4/PmpVnWE6AijeHzu3j3o8oYMTb1ogwTtJuqvEWWBwaA
/wJbr2zubfcZFMJgotDVbWlOP6/URAZ8IAZ6B4Xzii/3F1ItondG3b93SW0/5F3FnzoJJa2l2meK
6ecQKQXsTJlSvgofIqxMQRMfZk/dHhrn4n4/eACf6kcWwyhjYrBkw+9pHMYeW4ZNXUiRWY4a+KIY
E19nQl4jcgR5aVgqzHtt1v+ocXpzz2A3OGKvzWO7p81POgEsJ0BW5cMXnbZkF0FF28SDYaixUmKQ
QF13LQWDZDhU0nRVGxGE6FGsTFk0N4QQ5N6+LFjNJ+4SzqydyJ3WLOQkZZJIlPdfzn40u8bVGHRu
bO8eo95K5WsB82zLJd64f2+kao+nNmItgwJS3tWGMfjZCNUaiYWtHK0OJ8Qydnmlie/HsK2W7U0t
De3p5rPa0/gog3648W9oVIlUeLN8xS70PNHzouRu+tpuEhNPKYgehqz78vlZd9glsL/z1bRKP47X
HfrO0LwjfGGXJmoHM4gz3eftJdD5m/G9ANAd9/NoNFWwA1iBrxcMCYnWNQ2hXsFTmi+EgM/NlDlO
7ObOal1K6EPdsrim2JX6OpsfPKncB1/bZJnnlFfhn4liKdL0Ky4yZ37bVZ/w+yX2cchFAo+Cr3i7
zzbxNsyQY3Cn67dC5ZsLW0mEw0B2URlPcB0xTQHDBqkzb+2iu6lx9qcGGh5WLoWQO+0Rq7uRPP40
mRhx/dVV/WaMQvx/+HuInv9YwzTn+kxvybVQOume4Eb+1+jKWZiZPRi6seExoqmaQvcQBPmeeWqs
YaGfclhiDpitiG75PBtCvF9XeGmDvFmRtleli4HNig/KJTkmzQNRnvkUp6yYPMd8fceOArWTAu2E
ItP4oliOWU/MjzvK+ERTTll0UryhCK5fasPYfyqLS4NBvfn8Dk+nPO1MRNIIiS60NMxJi/GvGggY
8efzUfX8TBm0nMfg3ohYKTpBwZccXFzpJkfp3ytCuCHar561LpPIm7/73lIUonGzyXoh5FYJNa7f
Dy8qTS/UZRcLreEtxJtEJK4En0NKUCI5ARLVm/n2Z0vVa70jPB1nDjzubvviYmD5QXdOP4JrW12X
hBtqwXhNM8pr4zH3dMqKEJ7H2ISVe0uO9ts7yvWea2hj/AXum7qIn+P/dPPcO+LGHaN3F1TuBnHs
prl93qX+bJTcpeROhIA8pfUF2LTxVnEH7+xX2IirZf7TpBUxfXAndo0gyxftcbBTOIXmZYKQVpWJ
PARvD37WVzR4U3gOa7gl0NddvoMLG8WWRbsDX+72C/o+kSKe3kAqycvFQi24V3okCT5kdY4+/D3i
wk5euPJWcw3dfwgHip7t+24F2MhMXX4FgAFVFP2XC+X04MCXlg+1lT3GU411Lpe/fpLibrWjgFfq
lSBQ8jFEylm2olpe4jCf5f9JTzDX9mi6FM7SMKEiqLnasefFbyxqfmxhlLNh6GUI2b6yxs68EkAF
rpUT9khjXkcuMetNYPUEQ/IOyxpoBhL+cWVQBOeysCFwQiz6CLaxAh7ukkDoWdL5Vuj7aqpPxU7s
yyk+zYdAn2xOygFW62xlJrWNhZ3Nvo50Duaz2qYm6Mx9Kz02M6pi1oScbPYdZnRq+FUWfIFE5pN0
zsMJPL8g3oG88RtFaI9bVsmIL183V0/doT3RtvdQq0TvTeQ9tgCC/ClA40azQwFOK+e6eenQWc2O
8g21MVPABzMIe8Ql/zdL/oEgkHajNfcrWqtpQFI+W9WVJkeZVVlDUlGHC9RCRER5bCLITUX1WVAR
jAE+tYIv16LwYmvcDSfmKXA3HmqIB0prTdxsKbyxHSaIchj6EWnZBY1kGuBaBHxS1qD/rpkz9U3B
5JpAdoxZnh02EiqTozdgVLu38bNCEQ9yc27mTaI5zsOWdWrxkonBBnDb24CNea78b1rtOiLzdzvx
TtAkjQv/tVHQDM3ieMQ4UZ50HHkzQA8GPh30N36rzAJ5nUdA1tKW6CRIu1JlMgsFG7f/LCg0AHGn
aVNFLAkQCHvVjpy//5+XSGe7zx3T4I9B+UU6uke6VxSjhSh/aOI05erUWpfQ3wVT9TDLAAvKblce
Fr8Ng0CXxrN6Tb/oQtk0q4t83SgyINA4jbzRcxbHmCgn2dUvFSwSijf4SP3XHBGky3iJOaBJ9iAV
1cs42R/AnRbhJFQo4Ja9OKC009ygLCll1m3ze0lamFbVGGi+0munhXrkFwJEIfVtHiP2DnteT6Uj
d5yTik/0KWh3zik3rYcyldpK4ilC7MLcqbl761AuGmHYMQ7MS2r6ew72uANF6UzKQszjP2JrviX2
eFkhLpPT9+Sq37/BmRihSBQbiOTuV/V8aFrzQ6XXQgl55uGMuD06oekxczNJEVS+yiUkBs3ttnKA
b4GwpMrnzaWEWBPXWXeCb0nyIV4kbMdaeE9K7eZEhyaXj3sXiqEey48WNKTcYVybwaa4W532DaHv
nAGPXYljn417SgMXJYlpZySeA91GIH4BPhw+SeaiRI71K9kBqVohm0tjTNW86icBR88raWYZ8tn6
uPnFbH2gopaG4wFTdhNt52RV/6yIhSEl33sJJcKMR3NFFW5R872ejxnd0ML82Bo+lwQAFRybpou5
iKKywUxIg02kk6+/YqQ89o+0s8FWW7MuquaJ99PPq4ehc0QzGJRM/Ot6lD822vceo+mRs6qQ+k94
e3wTJwMmxuHLMajwY7EYh494BW4s+7ZKYYv2sxuiJD7sBDtLk/xkPi37ZHq8SpIrZ3/QV4yPBLvT
sRIMqx1Ru264ngaknVJMh4NizCJEQ3KB18darUFUsrVcFfQmyp7lbOPHYBXQK0O5XN1GgDux9Tq7
+0/ZU5QyImoE+3ihdH246yhUTg0JTwMAIg8r49iYdbo3bpw/Is5m8HUK5VTBwILTQvmpGkX0qTDJ
crIqq64Z6kBjPzCx/z96SiFViiBfw4ZGrLAAdgeUsLL2tHX5uA7AxlUmB2crk91+qkXdsTShXgrs
WrzNXnmKUkx2vjzjfEMz2+Lkn/oUzXu+N6OmkjHn08PKC1SzKRc4pyUuN68BwOMa33KTCYvlSSRy
bLk8EWZu/eus+Oab5E9U/urLCxgCTTW5EyvqUrNe8K0H5EvfR2hYGmjJtiNmD2nOg1KvCrRM3FMS
ak+iijavBVR3EsK8YRmNgLbpDht9Ytw6veYi352y9ZofGsf9ZdlUY7OVZKUtiHjS1SIwEoMMiops
rWauGvdVKra0eFDc8Qs+yJqWtQ82qj/6RnH5q+ZzI0du/G6e1ZzB8weVN36l1JiKckOqMKDX5M11
zylXVXqkPdkR217l4Gl1Y9+pb83hXBkp3Oyzzx/FsxKL/YrPg/ta+ntf9mv9Hd/QFiIR56sJKDW8
764MH2h/NcArwgz4vWrEsTxycp46CIJPimgAgMn7Bkw0P6n4CFKEcP1xokkrVVGQG6vFTg3EIgUe
FuhG8jdDP3R1YnVpAs4hBWhDYwb8MGnASfDEQoTGG9ihcZSDoU2C/bFNxmoEDISsLtYB9hKdb8tY
2ovhBJN23QNc5qn/AqPqQdPdtNbmWBoHOLdKy5ERwt992tBe86iJZPHoZB+57luf1BO2bNG6qhkf
DH+HjAUkCA0yVVIawb7qalrglBc5ffDGFAm2Ew8YhrihaqoizYMKHy53u/xWjYKhOGpJVKpwsFMb
6fziHbO1kpwEJPTjuUWVmhK75L8mb4Wz997zqptdDuSKUIGpmvENfh1/RuxustbZywui3LQZtLtz
VHlnGX35yRsU+0EF0sfTRk42GgRfGG1Riil2qTg5klI0Sc6CREwzB53kTBV6ivBVAsPKEM4mCIyh
8TkBM1MiwhttbCymQo1cCmhzCO45C3eCi0cCQ3SIV29778uq2hZYNDA7P3QSAg0KPkjAGmtVMwQf
XYbiLirZxInp/YwPU4e0qqF7LCTjP3jsCou8dWrFoR4JaowK8qn+4HIZuiaXPzJBD6RxacHsRFKV
bPBZKB/ytDkQBSAqUv+eRYBhTSx0JmGHdaeVsy0pS9yIA9ji1BFUFDqFMSRiJVfGFNTuR4lDRE2V
Xz5bAjyb4v/oQ6eg1Q85r1xPqESV60JHJhtkApnYcxtxSPvJKNSlN7SaJz7I9UebrCM72dsOW7Dx
bvthYMVKiJlTTZ3dDVFiMidMygP2sHdA4K0BdbX7i0+W9n66mHKC2ap0lWeIWXSQDG8VxxrXyc2m
laJXqdaEaEF2oC9WG2XI9t3A5zY1TWrUcVxXMoBkOBO2V4/in0t/084w2Tm8B406Fb1yCjIqTdmj
tDANIFKC7Kyv1umPBfFMJnsQC4B5R/PI3ZsoKgXNEYVpSgeyWWVEFJNpoU30YSoQ/8pinnphSSx/
joapYXIskqLVFo1IzfUKr/WLzS39joIGsaL6LB8PyqFcQT/JFbZ6s/UxyP26E0IH0bxGegz4QcFN
w7sTyRnuhziYL79TNweO6JOMk9PITthefSHmVZaByAOi2uoZJSrbNYCE0w6d30+wG5QRkBakUsEe
BSt0vTaiGqYBw4u1SkJbiMLaIarukvrAmjbeDwfDc0idAYVEbcxX7w5Sso0uKGy2wcmPvrTDjkpD
ubSQN0AELmkP5ydRfEz9UWC7RO8M1ewnITUEpXr4lZPbZ+AapdXQO29fwN3ijmy84tgjx4Zy0oQ7
h9B5dg6sdlYUqpQ2T2Etv9tXoFnY2KvcdT2/oA2BMDQui1Nm2aSb6n7YyzK18f2DyrUfusC5UJeS
hgylifBSwcNavRRxM4tQhTRGSrsGol82GjZnO5Dp7ZUP6OhnVE31+f55fcFgIXF+nbKbB3lhQ8NW
uh69nSk0NqE3L0FP9EMP12mQHqssdV83jQsy3o8lrnQJsMI2WnH227nVKWD/thhtiE/TkHYHGXEM
HBB9QdkXac9jFqzOlwvfNb1ScmCfjVXYX8+GrprdsjfmpfAeuQ02dguuw4GPNUfhi1BevApOihr3
aeA3kyaFuwTTHrTDwCitKWSuMfxZ0H/xv1tM41+bE2+gO1UIGZlFQiaiR/H9nZteymrhEauWonG1
93Hrhkv37R/Ot+300xV5usnsdBFpk/x3qSO6UA6bGl8dcyxMyJnXovN7vgqLk99LE3kPBj5uP/pe
QkDWtEc08lrUd0BnBpeuEE4BguDqO17A5EXOEV0LMi1hGS0+GBnyimuklrryYmvvGqXY97WnDe0k
QZ7WJatSTm7D2M68VVJmRm6FZMtBbqXUv73SupDNAWk4SN2VmpVzUUYb1a3V/b5eHXOOIs3omDpg
c9l6CucnJCq+kywiyXepQt1w1KWyXUGQwt4f7awSTqZ23O/RmyFbiOhbsTuSySRAjnZFhDX05mz7
SGg4FIV9ZLil2Q0/gvTHxerM368HKGpRPXZMlnAE4nIoBNRXHYuZ0l/1wbMwBdPk0SX3BUeXc5VP
i8N3v2B1FJUm18YQbcSYvsn9wZS8kR9B5cN7bMilfPCSB9IsOgVmv7Su/7P5FiSTZL8r6yW6mCqJ
K2w8KDzZ8fDYf9KzRGddGs3QKQ5UNN5JM0n1f93G7vHAVQ4rwf9s4EH4xNM9AeNM5U16nyMB1HoP
/zoQY1f1VuYoWMSg9c9bZoFbjWew2jB/QBy/zecrkyW0QsMRmM60du9GhO68b1ruhBAE6TshYbE/
9eXjz0fOraj1DlpFtkXyh0xnIpgvAFcWMGBa2Ox8QAEmaaHsYGqAAgCQ8EhP10td6M4/etDeftPs
C5842Zg6IqkfEoDs10zgBqRFRIlqic/JsPkcm8ClPL67bkZ3fWxgQbfeQwFAc3UdmI/bRUmdFnYc
KyFH27KWpr4Cl9wlPl8oh8RUZu7T7DXPLZ3l4udtKux1lb2NkyNXuXi5z0xJQbRjHSacSIgSPSZ+
MVCBdbKmDjNsNwwlyCt67wuheXFmhf8ehOUqqHpbYEaUo58HdLqSJo9ChDPaTysllCkZzXgl0FB1
pihbmagX+HGIjh6NuWGrDNztPMCaSlxAy0iABOp4exTxGBuIGkg3Mp1kAgSahwqRRf4mFS/aBMTn
ao/ynS1ZHDqF7cfAqQcNMwW+QIleUTz1Iqu+P5f7h+QHdtTzOKs6+DLulYRpGAOEHJYvzV6rzw/W
zPpORYshqr4YiEG6AB4D0V7KmQXeslfBIWzDLfzMsAhKQooUsR0+UjZkuzGOy45heB4eGoBFymVG
MJb5j1mqIFaBdrqzOIrs2BHXiLksePUCM8VNJJ9P14LiqgUwsCDL0WfkjSkWgf6flhj1gnC7paIY
cXR0J2HlkiFSTrdkgA5p7aC/Zf/FnOEwXQjAUiLohh2Qyx4syt3XakrNTQ7xSuJPjBqBOjl1jVvG
rBWTWxebFpUkK8lUB8MAakQHwOdOfbAdB3MkRRD9BE3euW1Ko2mHkB34eDjl0qllEdtQ2zPyfsH7
xk76++k4mNKLpo71sN3yX6k55jK7pwVM8zCVGkUKlpfFNPYuIZ68/86qQOz2vWk8Ir7vtnu71F+S
zyexixR38+WJAqKyDeW5+HFv59mipYxeu6iCci4UhL6C5SIr0KEeKxkwMMg9AtHUPE49kDcOydVE
ylXy7h7BOIXS2GCIYeeas49ej5DBepsoo7uRKGDzFfjIv1Mzx0JnO6y2ijYJyvGwpjiQIze5dtq1
dg7AugWXFQJCu82tqEew2MhMLEk/U+aNTFMYC0B1yYQwgHgjAu10OJkAsNmTQH9hyYIiijpyigUt
byhR2pMVyylX/0IZeM2bRlbEWnRfhnjO69Fyg6I5RZnev6XKtYEv2yx6RW3UAyi0zxVUXREE+EpF
ebYfgttnIddBR8N/R8zMeeIPyWNMVmAd+aWFB7EeGGxHWsKzhWZKpPMeFJRYqhkR39FK5K40o5Pq
8eIO77Pvfjsg18xmE3EIsNLYV5BMAes3oVTUy2lYYMaKyrRgL/4jRyWDwHjM0VAhYU0Tby9sAzl7
8UVtexFncbDWJ2tIiiHMWQTXzjgyGOoj+FrrFR1sCeVgyujjwzv0SXaXs+E9HJxDSknmllpnd6BG
R83Ngf7wZsempxF3v4sgOq6SaHIbSBXk47QCqeF+NZtJKvcKMp7XU+oPt1v51h/WmaluAKIAB+Lo
nbEfN9j1jaQRDNMUkdHp7HI4bx8LlxP8wNFJlbcKYC3fGhpXSHo9/jihQ/uhaWWEdF/9LRzyIFGN
BW7dFPgvzoTqfQ43RKmWcWOCgErSuoXtw7/iyUjFsQNFLzm9BXHQDiVdxo2CXjjQN+3gi6Wgjw9x
0m513ud+9TTELzsLAFm4DSKjC3LpZf92NSnKr/WfSEG+VJ6ee75IdPeUDOJJ6uN0snt5g/+EIDAG
o0FF2os5o4MknQ+01fU5JH6OJw2It32Duf/lMKZhwZYYha7Sc+wZF72FjBvL19CiVxh9ldNlSprT
M8omxB6QE0OD/V+H7pQdkdZcRFSbita23mfAbfQkh8n34qFwDxpDpHb6pReygspoDqFdbH7dP/vm
xoNfeCzlviYr1uMzmuMJRIMNVORtd3rrknupfi40Ms+7uFImERJuEm2kgB9/sL3P2CQZDzrRE8gh
G4XKLfU1d0k+RHO8PC/5V6dF6zN8+hnqjj7Fh96oD2RZsfuqlzenKhWRAPWrGQuQ/TFX6+4WkaVq
EsR5v2v68CbTrwS5YXjBN/j7SyYDFTKnAMNWwF09mYj8ENH7xfd4Ss0ctWKEDYaYTY31vhgj5hpq
3+mLN554x/2SpVKWAuffgKulz30yJkto6pwiSTd7qyHE7bp8QlLTfWAtIkjWSFxuF36ZHWkZG7Ik
1i4CvCXpVJ4DMeLkUShki9/SZ5mWFrdUVZ80Ael1vux/r61VKzWA1aSrSCgKL38pPxO9JPgy8qb8
8RFchn/VUhStMrVR80xmbEANXrYBSrQF3ddATqPa8t1mDU9v+pxRxCCmUcQnOEqHxgs5acUMY3wl
e01Y6gjiawpjIs7ZG5YTmZ1QgYCWk3TW6f7XvYOjqEJJFb2Mf1ht8sFhX1uzhgwBcrxLa1hskBDn
VuRGTHfzOU2rBRaOQCh5IanBShhJ0j7tSGJfNbJ7UwkWat7vPGxfKEclkhD797gwkLu8lCq6IbNW
X69S6fGjCk3B+x3Rr9y11TyEJPNnpD2t+H0XdxaBbzaJgVVcG1lVV8F3HYhM15qzGniCy8j1rZat
C/aket+H89u+zZ8nc/P3A0Ulm82oD4JH4ZS8xtBzQDjUPQbqhRQn5n5XN0EEAqaLVUzLTUjOCuIi
2zJxRq7iyEFhCFZCKW7UMVFOAtw3RjLcxsu39VxF3M51eHbHwkUOjtFyVzAtE49TkPYJgfosk4no
LUHBfwYSEnPd229n+Zyd+F4vBlvRFDYIP9GmCLonsqTM+lOc6AxxaLiJ9Jg3H3i4ZBjBq10Y8MHg
oCDWEBzviZwDShYXFqJu6kt8PrEU0GMCe4FtrDl1+KxN7YAZgKmKrp0+JDK9IbmeW4bgPv60T5s4
kOw3BpfX0fp3PzKT8tDo7ddxWUHS219uZSd71+PE17H9ZW1gQyO8y1jnqSH+sqLNPxUTyN7N1m4H
KvJhmn9IRbRA12ZSfTa3mt9MJE972j3oluIxWd2ferC3BhyvDjojZHDh+YbnLdmGy1EK1aa/MFxY
ZECtbCqPnsNwveut6PmzsFlagvuw1Kae+wNqAYRwwv635mPIeGjgKW7WcupatVo7oSLfa+5LBbyu
YvwIwPIL7uwoikBHQmZ4xyLODdZMX6D8g5UM2DfVspdbqwN/e2CV0k346XROYYi0A3O5c8LYleZU
ComcUMKlaoISu7Qym7/CLyByq8vY3wV1Phic15mfy7Y/B4piERuzHuFU+7UyGmKtPXfP2vmNoTUx
VAqk9mFPPXuMg2aJHuTcXo1sDB5hRcN76do8+33tG6Rcej6jjwDi+jJFgPqVxY7UH1WuTTn2l7tj
V2NBiIr5j+pmhvpfy7y+MZ4q3tmqpLYEOqTBCOAkABaeu6OSpIutL/+t31CYG1ZZUuaV+spZKW21
FoT98zrrOC/15/kjfakpuXM6KHp1AKTTuzwh+4lurQP+0qx1OTosUrAFVruXnNSp0DLjFT6vpKug
qWhn++KyyVkuKQ2+EH4mZOFitsqo5vynAxmbF5c1plCtqoeUsRiMtlIk0J2A0PlSagrbllogBYL8
qHVOj/P8vLNjz9yXJNCJblpUb52EW38F9C2Hu0WpEvv6eohctHo8firBPAmWHLqkBvGAwsbleLe7
c6Xxc7xExdmaVNaRyvBhyR6dVa5n9NF9KRo3086kou7pKhgcpRSYhCf2d/g/P3ozF0YDWMR4tFrJ
Va2+MPZw6AzjpwviobBD9i0PYHigc692FwC/iAHQILrSy0qTM8kEhJjWm8SzpO9WOUSVIAvkrXIR
gyB2GOMFclxAftJDfplJ2VAcZQXYqAiBlBF4+9HdJVZKypUawYpaeMi3VA5ydQZvf/RKOyQUji7b
DChM8DyCPfbeF6DXEbIrazkR7cqhzyzr1suh7AtDiX5BN00nbppuyzrI615k/rNGnhs6dEaR/A+j
tEBnfyLTbaXzPUGvpYncmkGVX5yp94nVc/HARFt/5AYF21aPvvJEGDVpVG1vYvR5DgBfEQBRop8n
fSKAsETRg3fDN7RJIV1oktXoJLzo8ky4NqB88qd5fwl35pqru99eqPTmacuNziksx0fp1bQ1KIT9
YmXCB6OL8FmbYvSvETe9uxkf6Ipz2R8hQWWezD9XAIW5clsesMWRHE7okl9Luju0NDKBE/xvaeVW
SzFYnVbIc+1EPKzejFWtSkE//k30YMN3OAYOKz0j/BSMSU8vHWIcVdOBgmHiSmzNf9siIFKo8h5t
7AvWTEq/BZYXBndM97d+WsfQlX5qN5NDJuEhVpVwfWtvQYsVgE4u3TX5/vz9WKa4tEqjQf+IBj/n
AzDJUuJ+w3WQJZaNRKMfzULzs+Ab13Izz6y1tSVmv4IpN06/eLhQjEZDy3UDxjHlmmXWVanTBsXi
YhbWFJbWot/TMYL8EFAmrDwE5ojJ13V6WTydva44GO1J31dy2pEbChBoqNJ/rOh6iUcKVK6ZGdA+
/ItFP7BYkj1wJcvTEKls9WPUqvDpC6TZJel0eb+pDFRNJbJlH5Ft9N5qXwhU6WHQVA+/BeJBGgKZ
YkAk/JAcY6janShdPH5J8nBtogehCZ111nVm2i+0CJ6On0/KVvraJYh5HjZqHJo2CoH9GyeON2TU
V0ClVhPU/zxXmeOiViicN9GAUDayWVMcYtIgDldlw8p9WoILP8xpSvE8LJa6MzY63UAxG17YPlLM
Z03BjNW0cB2ZBNJ+w8UvHunp1itUhZmR6n/tuoHbTW2ZWYUS2RG6grIlcCAdOCp2hfpL18k0Taud
Vuev0kegGQ71xTdChS5UFdeAQrv+L7cO/5+t6hvbPHH1aCFNu4vm9LoeQE7BqTZ3XfstY4qEa/vw
Az8nqQYIwSjhxiy0acT+b33a1/Z88pShuAjH9icDwvUY3i+d96EfDezrTjd8YAvdlAbNANFy/nSc
Vl6XW6vO1RrT7zVjNzD0+Qtjf5/W/LLNvfWUDSrNi/65kzCthxXZkVyfXNyt4hJgM873+BzJArGi
Xpjal+lpM9n/F9yAT/mo5MD/ytiVQqjy5y6URj7cts7wt3dEBU5nWaYBrlbuBOpsNTN3a80WFase
U6qllZaRo69/rmFjQA62FFXSwkfh6fx6m5ZFSMV5P5SFsgOSvt61xQVDzFPlwDcXVcfM/TGEBZZD
qq9kWhOt+ek6yFVDldAO9a5EijHts931CbBfZNFi6xAyA3xcXpD7VTVmdBYJRXaeKjsiVOgqV29A
hs50U+07CnwV8SjH8VfJRFTvnjJ6S24kaHRnO+BQVoUQc/kCMMiID58LsyOLXi6NvQ5bN9iG8ACA
14DPt/uJ0jUmRRjjHyTnMauhRX1vHNHwn1dyHG2mKZiUBpYyn/9AG8Cql8nyUsh6FYFwbfnWoQEt
Xdb2+/zQJo/zLsGWCzLVVRxo4hsBoX77bqXQQLrmSh+RgLMHOOtzrgLslDfH2rg3Aboh45rnaAao
Q10M6WqJyWg3i5xshDlJUiUTQq+lVdMNQruEPuQCGsIk1Zze6kGZX86eAYByTUZFeTVp2lOKqNma
aa/JkSz9YOCMHvxmrf1TC1F+3TNADuJ0OggBsjnt6xbm74Ivo2DHWOLVtEChRUMjwTbzshiTu2AJ
A367mAAi97GbPLucFnQ+BCw2CG8YfcLU50b/i+0PqsZg4K05wwhZfN95Mnzg88b1o3IH4+iM2cvI
/PAED9d8+QSQ/KzkX+ce6BGwgkeAV1tKZNpyFpeS1IzHnyS0IxIBoyhi70MaPhOk9c34w33NuTzQ
0KyMQ6if8bEwKqELTV8/WYWxZx/7PtIi0q4Fz0sMJaG3ef5YwBJFsb26sL2sEd4oqVSd3fm1B++a
0iw4cPuVGd/NkH9ysm6wkAXHmhRRGuOof0wOJZUqQlCksZt8NEnxqjs7owOB34KoddB9GO2/k5sU
pBZwg6VgdqhQSlnSGBSbLH7qm2HtXUcYzqF4NUcer74JQdy4an0/BZtmcwhS9Ovy9s+hxPU12AD3
CLLgGPftklJ0r5ZM14vyjaD9xF5gWUBDguJ8Rz1pTPJs1o2pUeCooT9rTQs7CzRGE9NDRdj7URVL
abci9IVNaTS44q2Uqz21+yOFPCQb4rlzY3++JS1uCsxze5mN0SrXLrgNXvZRWYHJVz5WgXmFRSoA
Dq4AiXV9QxGMJqs4OM6KQwRgnMEg7Qny3qSE5pQ4r8Z0OHEZOu3KkI8U6nSUJWNbnwcAQpPvUNyW
/QxvrbXfy0+9z57MHd8ztQM/30OTc8hywIa+xb2/ejKpEIxfBTr58t1joEBz9GXp9qTBcf9JqSY4
hiZcFEvb44fm8Ow8nihsAGa3FK0dX19aohYEgQVqJZY8PWkLqSFoSiWKnh0xeBbI0f3RJwgKuFG2
kECyKoR+XSy4sHMgTVh/J4LJQg0AhTGo99SvaaynUOT7JxWTCUqRJyJzxL1sZxdNP9XqsinSJTIc
sme2XQn3vrHObBHk90rUqRP05pNMxjn6wVPiVBY/JA7G/rQV4YcpgEsT+2cdhqGGvEGQZQQ9CoXJ
SsrQo0Ytojdguab+SEXRLZvlp8KMVfNmFU8AMILG7CGUSn7D6cOzWxU2JG4WRuGWE0t3tKo31sLa
xyIVzdR8HSUv80fm0FvMolP8y3wuKTappTJzhQE3agb04FX+KkxLToZtA1/SgIVWO+v6uu+7lXKH
TPVfW7FJa9ODyv/MGeb27RGBtEj99DlA+ik5MJ2wEiZilVeJzJrhXSUg+RnvQ8LPuuuqUSFkoth3
64TxEvFDgT07dZb6F2ZuE+KE3Tftx2gJIQeCOBXv4v7V5oL0NtkSKxMhUZdKGLUL+vPgee/2Zgr3
EIRKxSyTYtaTtjZbV2CRaoU3TajA2BR+dhnT9VBjPCr0lWIlUwAvvcmaveLlA2z4Sdy3YjL58Qrj
JSnAFGg3gYSrOwFXNEUn7fL5U9P0wc3oZampY/xc3UBwTJM0aINAjul6ibIdHYiYpxFQfBhmASsf
7tp/O89TjJKquuE10MutnCKUO5QfjSCyBxTw+z+trsHXcutHlvbH/2hpaJW3MEQFg5bDw82SRhGn
YsvEfkn1MU7IpB4VrqxB3qq5GQcS7evv/REjKMUAEnfz3oLdjbu73VfHzRlWFWkUl2WzN8gY0Ww5
lgow74haL7OkQ1N0J3WDZeveFORhbO1l5qyrUgHrgpYu5tIeRyllt27+BrRLo9DcEqLTXlSryREt
i558iO9GStuJIW89QoaAnAUqJMtlI8iwnL+Q7VSt/LbPBTl79E5M7NAN4OHqKkSCzdxgCRwSiHs1
KdFCjYQHlbpifi0GntvjJAkelwkwXYSWxYL6mthWS+2uKr7fZSZxJVW17xP7NYChUVxLmBZq5Ch6
O8Sx8stg9nYfNtchE5xSes63jPtPVHoJvvzkzZhGoV1ob35wtHGA8HplpvhGLfs8qoGDfOdvGESU
IFRT7h6PhkUjFskHc97i6ZwPmLYygs39VPxtZv3H7uSxWJzH5kQKgaWWhCeyS88gCpH2m1Q+SfvT
iS5Ivh15rBPzyPuT7eHR8p8lVh/JGBlDIQtPMhG8UrqoKUSGAoqePW4AAvDoLkVnTjFGZKvbZSoM
3bOJDJDAJl3+QIj/0fLeyqY9yStpM6zdcAflK73bouYQHG/XXozbENEx2etRAcdM4IQDAiJZQoPw
jmdXbi7/mFa9+nxSOrbDwdiS1xNbFhcYctMaJBtdIkPzeng4IHtAYbtwFpeNMf6H0xwctHdUawa1
/P08GZGxB7G8uS3bHQclerEk8Kq7QfjJcIoC4e80u1UQdf4tG0lmZEH8ksEpBjaM2TiRkc2+avC/
IzsNdn7opXWYPx1ILgnDss4c6QCs46es4DUgvMEcMeMBj0SZX/OaS3Cf/XUA59NLkyTOJ0TP5mTg
cjJ7JZQY3E9gCLNtNrBU4l/pk30pyVHPdsznyFJx2In72ATexmyPpLYYv0HcpLRtaF0OzamS1Haa
11QDw/I8iDfWrUKPBQmKkb/VqVuyTVT6jkT96bcsMHJF57H9oXhhoE9VveLW2smYTVe/VUutn4hD
IfpGIqnf496npIfITU9CBkNWi0M3ZIh1h11lBjXkJJdkSU7riyJuErzc1kA1Fbrb+QZFkOxNQYhj
QHG+V8mvi7SSGvmWirdhVuhymhxHJWii8+pSW3mk4okW5cPwqc4tP9n2QTGihXTTXUe03bd+6mNr
8wXn+HehU79IinoUYJT4bBjAyfDhaZaX3AJMFq54Krn3iLys3wJPP2T4wXREHjAEOeE2kWIICx/7
+FLnLF5LI6fVZxToNgHFKu3IhjiaSqSffeOrIgC54I4rDf1Dk1YaxpuNGLvGhhuu1w2zKkkZL4zq
x0xDpWn5GFxe0UyNGGjBrngSUbDD+IPhU1RLE5pbJXPfp8gisAIQho6EmJSF8B8oFUG0N3yWWnAA
mgiDTRQcoIg9HmboE7vPxZfqNwPf13ZtsFlDOlxnyLNFIbHOnfw43uZROTim//hTMt2647flfAzQ
9CaNRh/yXh4fQzw+QddkiAVfkc8Y3jDuBOO1gkT7W1qgodLTkBbgLYoAZniNOgE04DbXEIF1X3F/
reJoujPNeucSpEianP8Z05RjrCSvAJOiEEzEmmP/WBN07qd1r6HueP+X3mT735sYLgJ2uurJoMmt
w3cKYqbLce5Mo7XH0UOVjzRNLio6NsBTvmMFiFkrzkE2KUDSPJil81w8AbyiQV42NJs5aZXo7eP8
Pdj0p9MgCqd7QWY4U+2r/mTcx+P6IypiG1/1JguLZ5r0Ak6eok/KgC7PeYhrH9iVc550NN4AppU4
sm1LE/BBu5Oh8Y6b48zgnkrg7IfHbhq+RMNPPYQe/Z8+QLkWGbAc/+CzJ/aSFEkk9bHN2xzKtWPw
W2OK1RAQU+R8hptMvmi+PplnnjtRqd2tl58Zai7i6tyemXe9QJVvLh+du6sj4se2l0aIms4roPeB
1p40GvffWd8JWCvkGpYQyuSheiD+lJqKp/0KXCKj1xrWGYjVhAQCpkfQllJ67XDo2s8/CLhFhRQI
0XPeOtMsuytckcGxG0i0KBWFBDeddRtE2qVWd9sjwEDqXjbSJA52wDogVvf1B8XWJUzT8VqB08F0
DpRvRiWS0PTcVNxAvzPAs6Tuudi22npS78IW2e7tMA+8t1zTgM6z+NEhNg9L2EpGyB4Jt5KUETSE
eVr3NIgJVRBtJWoxijpOh9FYlKKCYScN2KAnvP6TYaNuV23DHDxAt9TCvFoPLzuA9EhmhClxiRvW
ogJ+8icEmB5ZXKmgEtDAq5yfjipQGrL4aJIuPN4+T6eQ06w+3AOrw3FnL+TDofRq8A+QymWD/e/T
bpYXUK3HMe4wGv24uFvlKdAONJ/k/vaZb8/87LLefzspZxPN7ebRKr2eqqNh9PrPPzy0spi4kF+q
+oYq0QYTOxsm+hFBAnUhzpIg0wURyEfRdlZk4f/dXHtnfE2Q1iQqr9yLQoB9kkyUE0/0WDEFiHeD
keryQtODEtO6uTvAgJbDqfhEkVqEfI55qSWlIb4WnakLyHIUuLjYWSbrzmT7ki7dRaVhSYBofTNN
61kol3iudiUsNXWWrWVeowLUeTtQJ5rH0Y4wh9DFrqisUaZ0B0Jp1MK127pQSIcHvBfrZk5DXt5E
MKxax7PXqa8Yk2ru/e8oW3l7aDgg24SrPeQ4Csn9X3gnVWx1HRA3GK9iuX7pqylJeyz/aVncs93g
NzC3ByMFkXsiZKw7076tDB4VdirGjDZkrHlNoUTdbC4kaC8UUXWSjuw+Rl5nSCfOZxQqshiy5r4d
E4vnvAM0Sgk1dkea5mboro1bDaZ+4klabFUejV2ndNwvEv56LdLWLOrajB8XEWyJydyoJLMMdAa6
ckzM7d/i9HO8VjgkSdYWbDZOa3lnWqBO59dfbkSOzajFFGFLkEyX21fzGb3OTuNh/T7qn5sZo2sg
apOSnNEj+I7jQw0hqeaPlY0T100D9HYcLMOqZQxSr9BEL/xY7rS5Cu2Ttcw3BK5h4ZvyascBiVBy
pPW7d8U1C/vhLd6jXBr9wieaa0i1oKrLzHKf4vZkj5Y8El0n02UTv9Wi82bkALSyOTGXRGGq+ZAs
LP8tqt7YElpnR0dWu+0Mj78cbSE/1D6DjOPdCd1Ctij/iUovk81ko9HJc0tvI9HKmaJn1Lg9Dgly
RsFQ0ffWp5hU4hDSHgHKWfXLO8Vr4AHLDAEz+5oJzZD8bCNqqSUqpCfPVOxcGP/HV73J3f2yvr8p
P9Po4fWS/3ekz8BhzSzp6EMuO3+OPTsbmORtMgvSWhBDZd7PML6JShuwiksM7TJGxiUSgD4euza4
4vZwimAm9XbhI63uLxEoqhS//MHY/KPMnJxNeoDh4VHTo+l/qlLgNlilmrdjyTsunjAxxsBtP3sH
4DxWDjgGndXtNnsaPY1vKObcl5L2lT4svZWdQ30UZEtQ60JmnvsGW2Zqlpuo7R8TUS5xFARNTMyw
Gdn/6OIhtLHh+n9URHbjjAxvxz4BE+BXsnykWPZ7Qmm9RWoKR/XcrSWa+Kr8kD5WQJsoB5VqEpyf
P83E7QMQQYb3ZEDI0cnl8+czXf6e6eI65Q45vwzzaBEYKIrhDzKPTiVloeN5pY32HA8gNwCQ6MdL
og83dQGnHaX7UEfn5JThU9nB0VOUJkp+4pNhrM0xg8Id8ycirfjCyTXkxB9S/rMekGqHCMp2uIwo
ZQ9v4H3UxjDmet4CIozMRTpDDLRvdfNLVXC3ynV81xR1wCE22Rbd+B01InON5S46Nh20RtHWzCvL
fXXkIr2radjQkQLe0XXDopkplazPeLifxnXrqZEzXb8dweziv8622GdcQMB/GB4fFVoRzOAR7S0c
VCoBItgNrILr90KEbvCSJY3wI3jUUIu+QkDg3BDZEzMKtbLSxjk1CSOPBtXDcZWS9TnqCX1htD/S
KYRkVshzYocV8uThbSDVEpYczJA943cvIXOFKIdnPAYlFsuFt+igeZX6C4fGxNJMGE6DwvZWwy0/
5eOnwZEk5tJ2z2i9UbsRfwDapg77HLQ9S6v9EdS8taaAy86bxyxngudRbMtKgB2+YGl22w/msbNl
lfmfvoLBbt6GxYTr+GlsVmdTAFEdRX2O09aOniFGed43ya4iRTandsH8Ir1yNBRyIdZaEy6pd+Wq
HV69T0pIdDSXk0Y5xgu2rdxUSV9IRpGR4eMwjAZwWJ25GWlVvRugNeEYUKWGkC9R9676dCgX+csV
D0q+r7TDowDScbeUgUneCxQXnjptzs9qgaxkrEv/bP3Df4JN9Grs0whZOPFVyMx18EveaYwePSsb
b60Of/b72rtrcs4yfcO42zLsQGKzymp+QQYDxnEJjHN503u+wTYW8JTxAmwx8aVHqk+wpAMhypnp
uXNRn6cLDQYrK4pTtIaUhhY/jA3CMySz2kNRV0R8kEW3qVLv4GvvgekljZpnpOmVvDbBsCvwaQ5F
4ySo0ex+Yn+A1uyp7dhMS/5cHsnPHSDUakjkD3Y6J+G9FQgx7WcX4LcrFFfnZ8CR1Qy9Vr4Cijs8
kKOYeuOL14sefPsq/MU4CKmQdjW5s7XU0kBnrjVW6NJLIWlVHFJHDfrvtfVoxfysdwOlLsHWq5gS
Qb3Bbxa3l3Zckxv3yRCyvaANZUGRLzp6PJPzjBnbjcKrI5kC+63OblO1vL/TSXaIDiOfbPDd9tm0
wMcG4V+HoRmkkvUgt13xx8CeOtqmuAkvZ1/UVHKJinG6TxgRjQnXl7fR/bZYcI7+zw/Nv3pHMboq
fAQCzcDzOYNcitqQbTzv+9kEvyODF2kOFIJGKIvgTaUJyfT/flwSfINOERslOuCL6Hkzlredw5MT
KHAhSKqBiOx3mEuYH/wsKK2d02XALHlgdjksxWXMuXjBalHeF8gHVx2P9G5hRcL/v4fQBZB8nBmg
WuRwxPw8wkf/fqys35PhQxzT7Vg+7kAkU2U6iAMZODA0LdFjadLd6OkR767HusqmL443xLg3qevX
dfBIFqeEgZxAdSfS64OITyqsuW/UE/wjkFXct29s6W0EQOXeKqMBrHWvZyqeaHUyPq6bDwek5ZcT
CRtx89Bs8p0m5M56WQLbg3Vv4frjnlRHV0ZjCTG4lkAtk08HAUp+kPhu62EzsbJGCVTvxLbEqDvH
VzcYnynPkuXjFMkuo3G3CbcyOpUi4Ds/tt0nzWFzQljoL/aY/u9aFPKKVHLd1r6VBYyAlnwPEcru
1oZhTYHb+bBtrUSNyGbyhZpmBlku/iS4sj02oMzLHa09Lt6TmSpmH21dL/KrSe5TJt0y6ghqovZi
9u0gqzYlx8Rlgia+AUrmVPBHz+4Ona2Uu/DJW/kBZG6QZ0Bk/ZWjF2oQcRcUA0Qg3Eumk3LbsYhj
PF7ZvQLpaTR1ppBkXJULoiLIMe4Aj4QPA/+4ucdTs//pcIJTk++BTZHZ5X/lpekAUk8g2lDlTp0s
7kURLeeIRsH8AohIdMMVYtPIbpHPGePOuyXiWvhb8XRN4uCZvW6CWbLifm7KMiEdgj5YS+4I2XH3
Z5yw/u4NALck3Pt0p8OU25uHULxx5GhFTn3z88SNH07dScb9Ca51a1ntQQJbtL3SA0kU00PZ9HgP
OYKtrTWsQ+NXsTzB1nA31h2gBxwEBaXnG0KhlEn+NLMvU1j3jKdP4zdWZTcf5VuM/jB3XbdWmajW
wRodpjam4Jf/YCYN1bq2BBDEcjQcwCgxYdhP6VOSKN2s3ZRMPWTB4wuf5OlLc1I64bbtCK8pPkSr
QLNFZ9xRE4Umznk08gqStsut3AXsxMA0wXV0CFxdZ9H13S1qkHJH5I1bqbf+KWgdnmXkjyqzqfKT
Bf3JIlL10imML7zDA1tofOnXKykPi0nvLCAp51S17aot5KU5p+oi1am3kxqtVA5xLUY5akO2d/q9
u7Hd1bw3h5fOYfZW+eOOla0gDWv+X6ox3YYITQiolpG17GumlOV307WL8yaSFe57ANBs9lA+LXIv
qSA8ZQVIwVwTs/C8Y/6jW4JtRpjNPKFm+I0+5WjtrdwH8BeFXQwtXK8GCBAZvZS37CLCzZCOLDq/
d54B3+dZ/aPUXuAjQ+/d0f+imAhgcR+7hmWwXBFDyQ6rEOJte3lzgoCssQKn2MhFqogHIAAQGTZh
7bRHXTKQGaiUtVS8sJTS7myz/PvhbIJDshxpbQEz/bW12azDZpTWvS5UVOatiUYzi5TrOPr/j+Oh
3PozR+xePmbigO50+YFfQ/vRkLj6UplQcGaBeV7syRmHU0cE2/wugYYrYg4fkqG54gda/ieFs+oL
7ytfWuwMiSDc8GRIpVuS4GpUTNjrV2RGPwFxj+Y/2a1E/REAPY+CuSwQQDaDIdvlICuHce+YyqQK
yks6uD43DxYQMkMb3JduhPKLDPzw0TyhzBy7e4wsvi16hRp+cWBAMebFbNbA1s6hqwrLjyr0DoZ1
hkFPdNH6GScCxfirEywH4fczLuobSWhiQ8eAh2M4T5gszGrqSEUUzZWcfZjNBgmkY1MLn7T5A1/3
Klpg9r3apeD24iP4qAfSzZjr7XG4Ns2eadEUu/cVU4iXB0l8ay273y297CzND8uWp6AiJnUQ9WNj
jPIOv0R+3F4Ka8c8Qi6EJOaCAoEAC9voL4WBl62BVfe2Iep06YBuQQO3CrqdqjFU1LfeoYW3EmfY
Xx8S5zA6S/uaCd/yObRm/f5xcLPsAvMHziewGSY1ISEPYfOCU5vN5hmdcfMc+sLj+Q2dKBqmPtv8
X1dW/Nh10D2t9dRqByOtOpx0hcO8z6Db7T3sdHiTS8NiZ9fIFGW1saXOs6iPgM6uJ5DC1Sbl63+X
anuwSj40Y2pNFilHGyx/x4Qay2wYw+98sqmZK+689dHFu+uJY+RWCtLAzW9lb6yv53itUnei66ts
SaiAtqhqyfyhc+omqGO31S+jptcPWpYREcaRpF194kslovUhsdoCzV0av5+UJrMA0Ehd6P1Cpwnx
YkxRVQ+N5HpGDd+LVzg3dSclOncXUekBIWidzhfsRbvoknSQYJdPJxFu3hSjubgM6/aZoDQAV94R
o0NXzVTPXgTrskR6VOBFBJZ/8zlxt3OMmsPgMdJzW6+EVqy6f3wGIbJS+BQOULH5YO8acS1JH37x
WsFqWwqqT5yh/fc05pQ5frHPP3EUzXgA+FOqq1zjDqOAYFYkuhmFUB3lQF/xtWKOT4r6MhIt52Wo
YKcmliLRHFwTsoB8fq8lIz2LeCZQG0SBEUsMUJ29ChTysex+0X4R5/hF2LZHbFunrJqsqrIadk9A
yQqi2ax5QbW9BZmnyWEkv9p5mZNFSRef6LQlVRbn94NszpYXRIskaogXuNVqezMopYiUpx8DmPkR
fBA+aDH3IsmLtKKXVzo8dEabnWh94Y00lhJ+Q4LyHa9osmZq9OPAhikRpLHDcxEZXKdwMkyTQltH
GAY0W2GDEYQa6sa41lXuR5TwiwA/NnNOKswdMp1LDVgiWWaEe0J5OD50DwUxNQQN/gpPYrzHtmwz
vZEtzenXl1MB3STXBXk7LGim2GrnaXr04NgoIZo6SMX2CHWZeMPsumV61bvACedPcmfdo+xBIjyh
NaAIO2deh7nHjv2MvgtZUXvz1ypfAfxig4qYOBufO0suM+f9IZla//8EhwyMjIip5SVFUXjdqP3u
Cmp1eMebjzrc2z0RhmYaRZNYEQS0HDqg8lbrgSFlCPOhiHhbVtCFnYOaf+3RnxJkL4WXiESr3W6P
2JfspoOT0ALbiJpoWF+wDj149OCBqUWxG4bi+v0rAsIa6S6AWeJtoCwujmpJpAqxChaz842syTeC
Uzi84/ckSo4EI0Nlh/ZEzVnNamXSroC7CRExFOsRhvPv4cimjCvxAy9vnjqgg0GysySY1OFAnFV0
g4Yyws76WcE3kBgbaGzD6p87Hg4Ro60j2huTNJMw1GYuGhZge+a3WbV9gFfmu7et4hxt5LbFcGMK
u1+jvZ3dJ7vJZ5cRmGrB5iNrmumrTXGiKSsUOomfkc9w+V4DlIiYBjIVJfkVGQwJJwAdK0X/Fexm
8QcyaIsQAPvuG1Nh1kDMTDVjPbMxAVmpWAPr7AZftcR2CmJ8G5S1lCI77VA+4lXeNTE8G6T81633
taF3jBJkUQx5buNO9oq5W+zXcTSUp3fTr2Uhgdz0rYLBh5QYU9YYqg68+38efnc94DR4I3NBgz+6
okNkBHEpuoy6UQyTmOb7oG9bhxD7ezqW6PLYetKyjFg8IYK63OJt7EsdfBImmJ7xNi2yQlYgti8U
CmVQwnruH9exWV9bgbaENAtRsc4fB8p0aWb5Rm6QnA09NUHDKWG+c7EQNZQjfU89F5S8JUNdIn/C
YH7cgSOzgEC4FVQvTW2Z2JF8DhYGNAHhdkaXbeAnF/zrbOY+DsQhB7o/Ruu/AafL5gxQ5GfELCjI
aZz7oC/d4/OOzkWWMtllULEZmN44lYu0RZ0eI3d91Udxi1BeSjMlaLGDftzdJC1PZA1IH6IAPPyq
cLXEfEqaLxapPYsHYx0DRBJyOWNFMH39jjMFTOE6RGtCF9256Nh7C9WNh9lfFM66jqtq3+fNNGB5
/NGeeYgIWqpRgIKdeIFB+RTEX0efUO1fNhuP59yowPIAJf/+hM7zFbsYJzShlJ5M+ncBPV333NGu
FSXucxgdqv+XeNOf+ErdCLJizICm0hd7ofK8QOJOS+/aFuJYFBmjooAaxbxpE3Np9vGbh1mohmau
y5oP+5Oz7Fu3afOjLo/ZD8+bmS4g4PBqGeQBx0N93QXdBd8w+6I0C07pF35bRPFWSkpYhwengUPj
YKqEdJX5TE3zKNQ8Jxst3Ueg7Hk2NNuWFNYeI0IXeeONpSWuNrnlRyJrdbIRlClZhAggb0Hj26Tg
FijjLdHPmSfL+b7FtNk7sxQ6TeRk4PseGJH7KutUi+cj2Zej0xzNgE7MEXayz+MVmnvmZtnaU6zO
6GtoPKQ21PynCwuo9OJEQ90XcV/H2juZw5W8gXIX/zyQaJsuXKjVUt+y7mdYhW7dRnaCdiQjnPUk
woCR4FTxiCJeNyEtsMM1X5ZFjx7WeHu/9x/iNk5xnOaEpfk33OYJP2sR6iQpIsetZ9Oug9uNHdps
Nt0FQNv1lc52U+q13rsf42aFwgGXZCfRKhdUYx+RKJvJtVp8sK63C4GrbKgP+F/+vC+E4AvS+gPH
Vb2DqvJKFg52wNE+YZMPspEoMPo3CN+7BDi1TuZmQLasHrZCqX+qiKTDGxqYNtpv0fFdy6arXlJc
eN5zr3w7n2pTUMF6YSwmbCPhMv5sxE7eEzTTu2lNiTp+iSa1PyzhcHLOoU+esNnocFoxegOwE26b
DTENXfrS2CB7KHSlZ0RmwY5NgpdITEzJos7Dw6aOmJu3QkX9EHNrATLZ6Rbzgt+RUJxBRJJ4s30/
6az4JCbzNkitiLOKeFmpvx4tQhky92wJH52q0Pm9B+lHRUW2VcbuBaok60x0jbZmWojmbzQ6x+H9
ZBDNzeb+5ylN9KlICIn1m6YfHwZpT0lw/YMrkcL+CJjWzqBs+QiXSDbBtWJ0sH1+Qf452qpPQpnq
gr7F4uXcU07VY+6jehlKJjeW0htUC448Ph7u2uI4KgelmcGQLUahQbVj621MF46rMkJ5hBLNuwxx
EmBMEclg5bqFat533qNnAmS5Q2HKpe6E9U9SyNcXsQ594yD2EzPIaX19UiToDqLpzQZ/eqzxQ2Ja
0nF+2uw6NASDFsxnOql5rkoSPmkb4d2y8yuzD2yfIpXBlLcu867E5WIAdco7IXGmkfGFTzDnu5uw
gYitIUdibM8O7SAmRiAmV5Pn9RklDSGXLruyw8WrYy8fIiIZ90HZHlwTfobn1On81P16EdL8G5yp
r9xj6QZKh7lmHu9GbKQ3Ed69CHxH+B3PQKP9eNR57qcXocz+Cte9wuitdZNc7t8x8nMGlh/BMaOZ
vCqo0WCc3BbHZk0iK4mqnTFuKcRV7II3LWkNTCX6SY4/jDhot2f6FZx2TB7vw3e7tfCaCnUZ7V8l
OAZwISDkzpIgFTjP7jeGQKGVeYTAumXTJXdoLMa3cyN/g77uFA2/DpghiCsShZYuVB2voQobKp+L
LpRD36rcMmvbHv86KaDIVORV/EPmxphvNNM2eNqtmZl4+2GrppRfJZaNC+lPyN6j3esPDzM4IGiX
JNSZYats0sd0BdgnZMLBL4v+d77H3Vz0hpC2kfR7iaPZD6Wt9QXQyApquG76GuenhAKO3ZuKEYEl
3PgoouFMezxFbrDANKE/RxHSoh1Kvlr6avf2Qret7qdrOu+XdHN+EI6E879jQoNLUJgz2Ym0z7JG
DQRXLPqhnAFlJgDEyMfs/o/7oKvjBIQx8ow75EeeLi57B5YREfRh+AK1TdyBCcW/JPjm7M5KKJOI
zCvkXJTZbSveUzNLsBRboNNMDqMkE3kODMF90QPapQ/2N4Jcae22oIWfwmA/XY9QqPjH0UIBl9Vh
yZYAYxSLt4cjRtXujcIf4MiZHfzISLmfM2lA0zi3Um/0i0u3nxV1enmao7hDxneGYzqSLLBxJo/r
w09F4fsBoQuqUOcn/VnROR8Mpn9OZ0ZhSwvoaQz1VrCFtmupxPjjMwdwyttHchTdFwNzNK7208Dc
wfR5UwLPy1phqzFULCNruNhJlO5U67esKCCBH4+1kuv3SfyAO1nzqwVgVkrvs+h+D0Rz2uXZDHmr
0ReC0Se+NxgHLuwJZerRqRLnl1i7bWzPuFjZdWoXiSSXo1xXlcpBZK1LVUIgzLAKxcjeOCWfBY58
ok9+Vwrac9s3NxRq1xy97jdYbS1/C2O81lYi89NvIJfp+wqIt/r900ixyWdWixdeM3I8IoH36DjI
hn/xlFynq5tRAu5wBnexrq0sdxB/lK5LSgAhDc1PfjzJhq/QPhkK7SzBbnf3W3cucy1PiJ5PlT1Z
4dD8nw==
`protect end_protected
