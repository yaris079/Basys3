`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Xof16aA8PZ/ZWd34fKY8ekcYPUNUNJRmKxz1JiSxaZqmBCt1WW8yCzwQR6HX9euSlCs9jWC9uyzH
fhjbwTmkSQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jKBsJ8VVQjh2HESzj+mJYbtHFXRK89kSwg8819NJRKYu+R40Fr32gykvrDTo1zoBlXc6wYLGCtX5
NWkdTvmHsyXbrKFePpos0NDg+dPe3ZVhvhLM97fHU6uw9i1V0wLQN27K/UHYFMriEOAMFEPk1eQ6
0TtC8SrkiAR1Xb/dWEM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CpdPeFEnoFGds0YrKDLyZXU9SjsH1dbuGiiYeMkYt2+l6dMijF/QnaosE0eeRUHVTLryRxgeY85Y
PimyPuyxyCwXDeAYTgHJKa9TNm1271437x+v5KCElo22QMNuW3vmWr4d2VXp6Quq4ZM5EWrcvNm+
CS89Sek709HhLuJA1LlZeR9/7gDmDHOb6/ynBQfkI5s7FFCpS5lFQGnx2greOZqwX+nXVaumzhWn
CcnDQBnAZIt1UCcSxbSoHexAbuozN6SerpXX4x8ncUeQPkC+enxex2XbH0dSpNOe5qgm6D/eHRXv
yLG6kO60Xcrbm6knJZ3kI7sOxNOUnmtSUOF38w==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KiZycy57VpEWmw/NRanBq2E3LOrVWqlG9K0bQZsZ2WJpL18eE5nZXArfKFcaX/MPOAi7fS5QUZ47
+hS6JC/SxGImJc/Mr94J/SJnapYnPCRdj5co9RBpDzl1FAIss7MVqDOxWUwwpt8I5YSbJfEVzwvB
9P6R0UVO/lZlo8jWADE=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pSoRFJqcyhOm6Urifm/M7yMn5+ru/yFuREroj1qvNcCcAjvY36hXa3DH5xZiz4j9J+HPUBrHLOHw
oHbzZim1Qnn8B35WbWZMuqICZ3cCHDP/xsGFYwCo2ErgfcUuCwOUHocCeGd+OJLIFZqjb0CtABMm
ThFPJGF5e5x6wT4sUlK96Igv2lZDnw0WPV8biTFPbWDMxhFoXFX9nEYxOoCfKip34Jo2u3OwAYRF
2r0kIPtRdbJr43N+ycl44BlE2+TGSapMSbKSlP4OxQIbpOg2O0SooM3toB4PtXMCh17zvBTx28jn
tgo+JgfP8WErhECH7N8gFzmyCAdxjk3BHgqLsw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40064)
`protect data_block
Ix5KEVt6NEHMFy4HslN/ldOCMxVYISBnbajTNvNtDDD0k6K9WIuY61FxxZ4I4J9DTHYEgOD7SHY2
+9cSih1IlGL3vPOl2iH6lu2KgVWdHM/Gbzdm+SmJaWfoISL3ctz10Mbdic3jKqHDEvGFU/EMP33i
t76p+1Y3LxLvE8M/zx60hXTBMfdPuwwsGp9B4xmnHR9EmiQ1gDEqm4zD8ToY7JOdA/MaFMwXMKso
M/bauQEu3rA48SBqMRoJJa3aTXfyopOjWHV+e2VFLpowBD3RCXPyEN7aX73PapI9/hRmiXNbWVqR
j9TvY3RV4DxZyeZdhMfasFCLBX/VTKZc5AJmGvWVORxV9CjJgJKiUnV8W/I/sQ0WaenQ43pNq/Kx
vDMx7RcZKXi3iiyjbymWtEHYgPfprmUZJy3Lg6Vdb6ncU1u8OWqxcKFZWOYeSqPPCqJJ+fJYlmBS
h6QzJzQBk9a1g3KfKrrTSWG5kaqe6LFo6AoTFUXGtc4AUwL8QlinurqRG1JBX8mCES/VRCXC0CJX
kdplff6YTEXCWb5FtfE0hLMziV8lvfMbHEP8Ubw2hs/IK2FAcC6aPtsoRUA9pASHYHkh3EYjcAUR
RPWFAC9xFbkPDr4lKX9vkpklVUNuD2uuXDvkMnTsHAziI/OZf8sWsbeCfkd3Z1oTCDWfflx4hWSS
KIdztoeewzHG764BgGoKHJJsbfuWJnUzzYHylGcrOzSErAjZzVUC2GpwdqUe18bort+KWUAlfCXi
zI1MJ8OymbvLn9Y7AqV48qz286/E8OUt+AX1rLG4DpgVbfvon3Ct/ZKsLa5WrsCYcwmhYalbpdUb
4DOYdxzlH3nLoifIJbRCRdHZ/dS7WMR7l4MDeFvYsgKeXmzUjt5vPBcJjhBEOEilnZxzM56C65cZ
GZRxlWlhPqTAxDuw8Wl1SH7eSIExt/9edfCdQONTpgNFN5WnaZFwW/w0CGV7uRlRweQEI8NaDLK1
OikVSENRKGIXHgqDfwVSsGFGzoU/9PsaRixwQcGBC5e2u1FDYpDZplQOLVGeFXPRBR+wq8zJIw76
Ur78v8f5tPwoGulIGQLkj2I/dJr4fCLqH8811DK0zOmTBrfTkzRUI2QbUD6TpsP1WSqwmWYeKYsz
gDwAUu+N1cEh2JBQfg7CJsAEXzeoUAf1GbR6npln4LMO6HNCs7WuIiS+VHyKKD4zfecSlvf6wM7v
bCrcql/IU9CgSVINSwcmOzQbfCimOzlWIikxHavshXkhOSrlpFMkc8cDq1GOlCPU3B5wXmBXZ341
YLx1CRnIZ+DtVFwQX5oz9ZRE0TH38vg/hxIriq46HpnISPuwXvPC9YgBDRXXxfiHXHIaSucckhdR
bGOfncR8n2rSyshIUTBkNIo3TwrkWO+4D6uF0s29zwM474i6lj7SgjQ2DpWbInF+gPI4xOBp1OWy
n+sw+RdEC2NeqkWtJeq7RDv6TVO4WtboUzUURIoF6H42RR5mLLVIInHSP6xSpxipPBtUyN8NOrPy
ojL6fmkp/7/xK4z60K+Po9i6mbLkjiUzwLREowVXYWD9oYpi92kejuofxmH9LG47oHFtI3a4pDfQ
6qjinTENfm4SCSPJtUQc6t7fZhQJg5EQiQbSN4viq1S6tIpTzd2zk2aoeaqsr2pBLrVcxueA3V2G
OkyoQs5FpByORoQc/tPOqxNpj/JrRSxgA9Wof/fRrh75SzQgo0+6BxVBKyhXaL4z9uX2ajcV4Mgl
Gql3N5/f8O1AfGvSB2rzlxXU/gGwqxl0aUY2Ac85blJ7XPf8c+QZC0aIrR0cR6g9vt2/RziRa/dW
SYnnY0josdLNBqx/chGsmFk4d6RGT6zRqpCfUG0aeV0vuruQoP6czewktrylXQFySJBMU1WzQaU9
LSkg7Hcw20HSlMxoNtiByDVq6rdjued6tUKDU6+0kxRYL0absVSkTOYjjiGwiNHymN1Zi7vw+oOv
RMudKp3XxD5DpxiShdGj2/MPdlv6wXa47zQf/Daq8D1a66lqW602h7XycX2Y+eHl+GqRweinf5X+
UA4MskCb8B2WtypEhw4HYSrIe3g6JZwCUdZ858TIsBSdfOScSoXZevvMTMEmr70/x0RxRc6FHupN
YUsBNewhyjU1UfFNV1tpqMkLLSDAGOMBLpdgp6AMejyeuJji2foy+TpQjwlYVbPksieINQzHAEop
65uQ80YJ+HUiDxVr3zQMhlDg+2OSoQN3zNa48bYAiHwiskkIyrYnJfHgFNtlSP01ecX/yF+SupZN
mT1/V6nb+ucvsorTVt03qZOl6vnTSP5n36bXhc06jPyFNOvUMg1qqusLC6In0//KnqayTh+fz4w6
DSDqo7jz4naMyFOIWR0T8PYjwJpOBUEeqeYm9hS8U+49mCaZsuubf6Bh0lhGcUTP8RDqzm0+00Gm
DndVEFrR0nnMgMusHkOvLytyT4dXDFAHAi5kib7YJelF1xu+DvWzM9Hl8oEwMx6nNMmh4YT3BCBL
ovxsDBGgB/vgGmagFeuRyejkibBPHGpKmMshlbixIrWHC60nnrp3QNxDvT4S5c1H+CojpUC76PKI
aSbcg6EnHU0o2pcrnFmtOqkryJTajT0cgtiaL11zVrwV7mDd3McVcvDYK1JG2GIAFq0Glhf7drSP
lhfCjYi6QeEPy4WKDVYF2ZldRTJjlncnAnqdEC3UG2dTVhZMLtBgavz9dMS1JcU3NvMOifPRcDig
+Y7w7hLZp9242X9WZZIy0CNM+kqE5CudD1SOfi9kngNR0+1MJ6HVRwXDIe8tG8Ywsroh7+RXRnnp
VB9MUyFTktYNDKrZvdO7hvTG+N8QFKFNs9tjlQhgNKZuga7ywFRO1hicdsREX6a/YT2R6xJV2qOT
sgVBs5t1ACmH8i32hBETVkSCqFetE5eIy9fyuI1DMYLCO1wvSQlpFTTWJKM+bhKszR+kDRK8EnF9
hlFXe0RsP+4VocrN68pJuCHIADtoNFKjTNLhbFZtO3RTC58xXV3WWsrKZnkLsTcunWes2NjrgqTF
xW094+Zv7Fox12yguLcLhRA5C6bxRgH70dGcEGwWJydkm/9XAIszq+o5DYgJIIGkF9u3WSxN5MS3
p7MkQWBJbQF5D4+DKgTBvYWD8kCGbP3apaQ39xFs4SzXOT1AlE7HzoDRGqSyazfqv6jcjg098pDF
u1WJ+dggJ6duLSSmtxrtCoess0qGcNDHllRs5wzn/rNMoE3REF06GBZDB97vRPPhMQWH4qG37dDU
nKhVtqEkNBdM7cFH4K8OpRztlZ3dQU/Wc2gDrHwOudDECTrvAGlm2VhTM25XmpPmicEjG96pgn7L
GqGpfvAA7a9/GID19A+VxJ6ZMd9UUWMpoWToT0Li4T72UPonQ/uMpUZjP+ep6NhGsGI988TOUyGc
fh+jqCssgc1J9zocuuMSannDejxmeJYZ1woqMsCitzLy5vLDlmRYcQtIPPLN/UJz4ZU47wr6F/PW
3Q4ZvzSl6z828TDiyrq1+0lPnFv+IHUY+NwOlikZWZQK9wAtlDYSPnfHbkMUhaVEj3ISDx3y063s
YxzX7oo5K7Ew35Sx5yL9tndRd5gAbTl0NWS5XFVGghN9qvZKx2e53gfN5EkcsiSHAmX9Sl9VG5wq
dMYWGrnMbgCe3NLIDBerpnQn1ECaxhDlbXwnJJINVYIcFO+pTGPFFOUYBjfd6SuoZO+Fk1JEEbEj
grdvnQCho0s6DmMae6l1XEYB5wqZ/Whhxg8sg5z/k/ZPUoeKvAvNLpM4uU2Gn+ceCQrQfBiiICSd
V9tIHWQjBfY19KkhQCcCZ5F+L0Tnr5ocezEahPC6Xbq5fYumsMkMTIUKmibUmtg+37AnqJMs3pmc
5tHuTvAbiyAseVPl60HUHYhjSjRwNGf1QLY7/KP9g2tCTKzjKqn11XTlhtyas57BDtU8LIMCmgOB
oo+Z28eK3ZApId1fIm7QdMEXbhW1wM6UkZFRke2t9M3o/IMCB2mpe583OyUr2UNU73Hf9norWV9x
uwp+6IVTsEJ+27+RJpmL0iozWdAR31qQpGmznOv6jXT8HF7Z06pLuKvMGgGBd+OwRrmU4nmzagPj
fD1R4LwhGV8qFcKdW/BGXZiLjaskf+bEOztJIEtjyXdSAWN+GZTKpfXZwDrY1MiYlzM6YXkWMhpB
wOUXG+bJu+/6CmngGXi/UDHs62uAKrcaPsFPkowbRjE5tZDvR28C5WBK2UVZmsQwvfw5VorBTmA7
+/qavL5JRSq528p1DeEh1i7ZClIZD4jAx3WnVjccF20UTKouq43WKugeSiLAH+mrcYtNAJzVSWmO
+vV58eoeDVQ0O2+t35I2GbywN6mh//s0z4Qko6SI/l6vU1XXxerwrCo8eHPR1qI8H2hkrq3Oremz
F+h7RvUmx7Rc5OLAc/EQYTBaeOFmSs7/+HLPHyNTJyp8LrIDHEoDM0KCyt5FPEhQYDn5kMhIdDNC
fPZxELcHdVL2OYygoX6FFvSEV0cSFD97pSjWSPla2riJtzsYxVfsWKx1xI/9SeICdKY7IA529UnK
n1PY0FZ5sZNphihtr6xgtrM4BZ4biHHKxhFMWmMsw8NcYT51EojQEW6BWz4uxisAuRmCb/ac10RF
W3fucRNKNu4POkZyaDA7zm91B3j9DgaYaw1Jkz/zhV7+NJ3qOfK2LvnWSRD0ptY8YwO0VwGQuMgK
z2GNL0ti0skXbKwMroc3EJftiltL2u0azSUNc+rgHe2Y6cyDgdzqulchM/DgiRPmvES/g5pBdNPY
kKKloc6U2wSt4ZB6wkaoQhAOtITk5gGgEEq6wk+niUyWtA0N9uRDy7jF4/pTuMbDvV5t5Jv9iqc/
2eusYhboPid8+YuHnBFgIA/FeIPVmjTgx4+7Cnfjd9bz2Vn0gyNTfYW+MVhNR+1yvHq+IeJhvNKT
DzURejvoiMflbTAH/Pv+Oo/yyJhI3q1T2SGrprlsS0A+oX7AMnzRINi03q+2x93n1GZfCJfVkAjM
0uHz7x55JpTAeRp7PS30Jran58MBPB+smMh3FXKvFYzBJnPFZz92jZl4CjjeIq/RFRjpwUzJx1u3
uPYoUfa5BZqlpDI0zCyMBBnj5NQzP+fKZGJcT063oIu2OOsP5AZ9AavFWgwjgfYU1I6IwzSsQtzi
V/7PYpidOPpC2MOCXugtGOvyWAJ1RkCTx+0VoBqSSzi4MbUnEdh1SWvlbwqFzf1R2hb8cPKTMQDc
FfjRW7qXug7VgcUFUo8Ew1NkwoMxm1WY1qPpbbMuqmoZMFTlFO+mX5Bx3+bwFg+hpmALMbPji+25
lotRr/jEGeMQF9hYZEgbyHx+w0yQVwbtkbhzC/iyXyRViXkVKCXNPucjwxJj0zlft63AgNscOsVN
YD1FqrViSyQ+iH7UqNoytZBiuo/PGBzi1tycFBqAPfmzEzMBi65MJARpI/RQY+qsRpSmhIyICauk
h5DTTYZafCFDWel1ndtf7UzTP0jjawby9r2h16PewVlhvARg6GbYIp134A1ch3bY7gyzev8b7Wa0
OhObyFOqFQcviBSVU2RXzW87AVbWQ4BByQjsk1Ln8HZ2wCSGS38wPg+wClqKVU8PDM1UtMuIDn3q
Ey27I7dxz47Ugd5JwTBYkTslIFaDLbhfcwtxTyPJi1Ojmkx2cGUzLt7DPAhK2QPpvNnQGWQbXAji
/xWsf+FE7vvv4KWO2Uu6X+3PtkfFM8oIpuH3TlD3TgGgQI4E8DDDJGYnwxr5gkeqyCULySXC4E6J
Had77372GjEUdJl2llJqh1ii9k1TzU0h2fdQ0EtafrBQtQFh2EkUVqCLgE2LSaQRQ5tN5Mr0XTw9
yJQm7iOCoWk0KAbnOqYLzh3A0WHVxyX2dYEmE5gJ45UvtjgCsCQASzquKzsCfy0XM8V3I8gCHcSe
JD6sgppKmtwhby77/GWEjyXtb3bdJzNwboDO+19/ZNtevCozIjSAq2UYIKIGbpajjd+GuAWVx6iL
T1J+iip8jZ7UpjkEBrWNJIknzedRg6pUboz2D5BceRRSyNK8rztFKYWwCstJT4YCmqw6EfKkWRM9
tnazFh6G92rF/rgLIxi3P8jLIXny3iZK/6CEL+9NcsndW/9DXSJ17rflvDHBPVhR6cnYWVXUy69q
7wbZCSOVKVvcwesEX1LDjLsNoPEdRmAoRr+wNUQ+AlfLoXfrAra+XZ/H0m5A1rtM1u735INCYcJX
kCk2tstVh4VdpDcM/tO203gKuIHhco3HswAXsCLX0wfqWr7zULGNIq866mLlZ1AgNBHEpMGLG5DK
E/1Vboq3cUmHzrDoS0m/jMMwnpK813ucESDxx+X2sXNnTr0BjAv+9fcDSM11ANNObSSjbDL3vv3E
/41C8lnDVeuxZBXKrSYo9ZzjfsUYBfCtg/MZffFHqgbZUKsXi9ft8PgZCwAQjmHu7LyDShr+7nSN
OHG1CM2cMlL3j7OtWKqV9avw6M+NkzHF/sMocFE0nsT6Qyj97qnQLu5SB7DDoEwIISn83+r36PCA
NIunSN1QjbJsThVA1kl7ezltoohmYlQQeH7QB4Hj0U49p8yl8eRL0Ho0iQD/ORsH1UMyjWzzJt8y
+URAVgT9Lir2CzDxvEozkQjmD62nAXGrhbndZAAKeaTID029arkz876uQNhFAdaPTVRW0VJHXDa2
znlfJExnkb98GuTQQfRbQN0WrQMWtxlPfd8XbA+i+FFEnfWH2tZ98X0KVs6bg/ATTuy7yIrVIXqd
BabatwztG7NwW/aBNqRYOxViLTbfHaTYXx4qeXZCbJYxmL+1wZN+dJbtGN9vPXwQNSGIFzFNO8j2
StSH4CbKswHbAfd47jKpPkxjK/NVutc6c216zhgHvdhnToZtDgCtVCcCBwxtvEqJ2e/mWee+XxpI
+iMPPXmSH7EMH/zrQVZzbrJoTtOC2g4/7VjS7VNdRuTk6httguBsJmu36fJ2WrgPHKGLYiHRoLli
dT11CXs+JZiJdd6Xdqutq0L0N7tgZAHgSivmpUfLcSnAe9KxcvEQQ7d1MLb4rlAUjv+KsTzsEgBN
GbuaVG4Bs9L5VscKES7lKURvPajere2sRzfJc1NteaTTj+qP8cIfQ3kZDWCa2+rJEiS9S57z+u18
PNOFiuAeQBn8GX+gaYv6hcvN26dj9aMk1IpO7Gt4hQ5DziytVUfXHj7XJlhLH9AfUZGDA0T+c/k4
ZZU5s7XpPVY/qFHViyCDuJLA2TXWE2mL2zRFe5vLQbdSEeRRvKQ0UBhQmYpWO6LxhRSOdEmpDoqg
UfSL9u4EMgaGNCPxtLJGpXEaIgwoC1CEssSXuFd2rH6+HJZnRDNOR15DhVBoeopwVCBvY0gyE4m3
J5T5jsU1V25HQjcbYNPzL3bI4EdE9GKOWkA7w3sAuHmJpAOtDBchM+NhhqOaS+MrUNH2Fybaaw3y
iO+cxpF2NUrrbIYeuCmTe+f9+89KiaogIWI109wznLsBWQFr1lojV4Lns3hoyaJBsCArF0HN6ZgQ
Z+R6TMZbZUOxDVN96rfYl9iy3L7kG/ESAnLHpmAZKPitkBDIRCrdmU3fkvqiueFEZ4z0YwKsLaQh
h2wCP0TaEdCMcZVk8kHoAa1kbeeuHaWUBlZifkIOjg5xwvebuTdZZYCP7/sIRPBpRM96U/90hkx2
2g8wikBz+6V3zpejLiBUPoXKYz+513yuyNpt9QHGNbCZUEnRVD9MQ1FGEqp88nmwkzE334sm/UJk
HlSfKs9ZZV5JJByA/4ChHV+shRZp5vmLT0m6C3zlUuAyWxj+kz34ARaXfS3ga2YKoEIV6jrid6Dh
SH0S1eSNvjQIOscOY0GFuuVE32OvdMP2wQIMIiLGh5DU3PaVSz2/4B7dw6P6ph9J2Su7kareGmPj
/3Vqq+G7VKwdCrSm9ofnpgBmvgjme3g/2DSr9LB9c1aWqEJZupQv5cWOV7JsAB3xOEjF640WpVsi
VY2vRiElLwOsp+8yA6tK+UDjzVfX/vCtHZsBtq9IQTnoxyu+aVDvv4l5TV3BalT1UBw69Lu5xAE0
zIJGsTBIFp8r5CsLVUDrc1oG6sIK/1KkKm5YBo8P3MpCyxcEHyOxWb9P+Yu2KXkROtE5OdOXttNB
jAx8cAlLQsltkQcr4UVHytSRnH2bjgSsi9RBTqJSBtNbj5b6OSgP2s9kux/jqTW4FEJgd+NsRNJA
HejMhAkRRR1NSfBiQ2xvAHjUfxj5eyJODeql6YxpjBKqjDFUmFY/X0Bc/7Le6QTCt26BSOLGc6AX
fjhrPP6NafwCfPJqxt7wRCgwX+0UaQRSarNKvh5qGqqhpTs8uFi58f6zmzdi+DwQvKu1cW4jiRYv
1LhUjDAzzhxfn+zw59ATu06xy1idyUXhFctAq698zIFBLiAB6caJJ4VKE4/GrvIa1/Hba74YO0pn
fKNG3oleS+l+yWM5kGw8WqmQ4b7p6q8Kdb8ZuBNLih0cwHt7ZFOfm5W95KZUvy/ydzJs3CVxzLpC
hlBk9bfZ3LLmLJwmaeG0K/go9LHL5KLLly9I0AQlIu72JMHoUFwXlG2eKKr3d6cyFm+IDRu8wOZw
ME4bnEiqIJQGVSPGkTySXSSwcD+6LGrSCmGt6t6PlNgc8V2nAuk94v/MsuNgWSiqp4Ad8SVTUx1B
ATD0YZhcqRYaHu/Z98wUArnmER6QJ9Bmiq1JDxq52HrXeCKMxtbtf4BL4w4YTlFLrU4b77kcfb7P
ro5HvGhG4qpBsUaBqJM3ptv5xOYs/2cMH670e5BGL2/Gpe7JQD4E6FSSH9yrZC/qTcYlucDpF4n3
B8qI8bg2vUJWPcpbIT+0lLWUJ+jp93owoSa7oF2wtliDbDNv7GG4JRSFjcb4gfwwpUjwWO2b1s6X
9gjtrDMDzoAC4ssQD9RSq9MXB6oMefsNvMSbkpdQ0j66pVKbaEdLEA4RMukbyrGrOE3kouHJgtZE
YrX8iqnGDd1fsInm5c+E3SvTg8Tk6mZDSwfd0mIOY/0Sj+ubBJ8fYX8Vmctz6wYHiZeOmb/kBfgt
p2ifsN4DHr9NF3IM+fyrAZILS4wTM1FMlJFMZejukSGsHmIhpO++VUfp/q6lMaFJmmRfZ0DIk4jJ
8p5cX8Xu5GQN1NmDMgRMNnnmSLqMZHc2wKy7fZV1kEV+4XVySejc1ZgAZfOxRldAwylzV5HFLEmA
kdWWhV284FVAJB5tTAVZS/H+NPmCNDKGnV24WinM36OA7bHzcx7ub6vFaUhrPJpGXK8rl9GWJ/rC
RE4hX98QDu3eenArnHrZyE+a4sMZgpsMJ4uo+Y2kUGOCHq2NXKAO726CKRqshHO31muChcI/PGoy
ca61UFsY0YCuI3jqgLn4H6UVKfZomKFhMUBdjFTp1itU4xJfrV4vdnpUN50avUIDdFUo2JJPBiFU
CWhKJBH9RqvW7wzFgnUHk4u7IltpfjBTa1Vhduus86RVwpYAH765MedTRnXNYY3jtjag74RX4r4i
Ol2s0g5QXqV70bwpYz1QHY4BjN68mQeZ+gKH/azQ9rVoXZclnAFR8sOh00Ysolc5uV2/opWksSvv
yWAcwrggAEvq1CGJAneIpwza48adpma/GE+vnVcz0dPznczDbYe2HlsPNEjeXFyDgeL62al+RgUM
XSRpvS6jza9EWYYGeQaM3SnOlx3JCze1ZuLXD8/cQMotjiH+ZcNsqBTR+JQqizGh5mmcCZIe1onv
ZIlDegYlXs+WKeVd8PqUJIs9n4xtJRxBGJ2KK+0Uj0o+/vc/ZEBKymW8WwuH+Ir956ZFVrAAqfRf
EMrE7ziyB/LS3Whp9+7FcKA8k7GW8znrNBJR5lP/Cunkd9iq54BhoHIg6+UYvkhvEppKM1mPecm/
BwdBBx+d5SrQwQ+d4DdWSQJTglar6gzPwF4F4mgCxVEJaL7AsgFJxC/4zQ1ulDP2uJoPS3ANfFQL
luk48o/NYzGRa07I4BkcJPfJLM2UqkAJ5UZ6Da99qrCTTheUJAShI4cgqDWyGGW9DiijDoYmnmyb
Z048YDjmFsRewN65S7jR7pS3x4/n0GaSJ8Z1qy/JJ+/NB4p95MVdJD9I5YF7JlnSb1mg1g7B3Ahu
9W/ZUP+jodhIZgrNRvby156x4NqDLPVc6FKPeuw2BogxI/UYGSSy7fkg+iL+EYy1GX9wsceREswS
FSd+laZXTMqD5b7DP4iotHpT8BQ89BjV9JnYtVvWnO2rkL9lHewb3QdRuKItpwfJWXhCf2FkYNge
tC3U9DjyPjjmdLS0uBNCUu+tzM8STy0Xm5eSwJ6N+g4kmzkTuaEH54wh2uzeDGNktAwqa554EyA4
j3sDC1K69YpeJdNfJ38mvEvCFC5WTO9Zu6WKrs/fBkp5Lg+oFbVFiUp6g8l2cqV8b48ct8jNtOx+
ZDZo6fseJltYVZmX2YIKqd1ID6nprsBVbHgAcKpwSNFIw1ec+FPJZvho8RCn8cYFcCuZxek2ZwZ0
x0YHkOfWQPnJR4+fQSFOAiMlSdnZQJIaLEqE6pPzMPor2HO2c/u2y5qmrK4spGI3sas6gCyXWHNc
TGQdtJx2djDemjY5SPsj9EN3KDRRLY5XLnytLKcgJ0ojZjtd/iLZOhfgk0GghJnKpzcHc42jgkr+
zEmz0vST4AgQppQeXrbUU/2HoyeXez+rCz/d32XsqdPl/te8sq21dR0YgJ+cs6tWr3pKTTJ3Z9ev
ByimJEoJAU/YlxnA8ilBIumafEK4jAOnVDau5jo3AxripC4O2YsRjED3KCHZK59JX3zPP3FonlhX
ozuLIbUrf7501FDSJEh90W9O+MT/fvGRiMIoF/wMWHGisO9q09iILfI7TJ5UiX3Ga2rm2hGBjsHh
ID1qxCdarLo3/3ZtPsAhbrmlknd/xnleEys+5LR0UmaSENdVjSzG/c1XgH8tCRtIHfuin1UTE/+1
A/wl/IfdXopIhaXD9Y6noSaW+2JHA4u4mQhdLATFEU9H48nDaDitwAm1BhEyHwF5oVFfATMBLr77
PXSgNc6+6rGU0x8sjNOlWzbFFFWnRQsIhqEoDVG1sULTDkNIvFoWItiiUyIJmpWaXYXh3ywyjk9a
Q4he0kCBC45j7V1KQBZ0/V/itCozFOfy/lhFAEhlDNfLA+Y3hTHEQN5E7hBrfbhLu497g8fHC/10
i1lrawnzhmmJoKh9d0EdeHeBbwKsXxpreB9H9yw9CHK3WwjC2py9F/zcPuu1HpzAnAK7IufT1ksp
S1tX1S3OZmMhl99pqZzWmjjMvwyfqTlBGYWZR6kpPGfcP6Czs3avCFQNYOBeE/PkPYjcNODyYDLk
V0qcAppUXmOn2B+Ckfm4imWZ2n7mPLzw7aYGsXDoHBQbG2x49PuRIgP9fQgj4m4o5dhVtMCbrtCk
scvs/CWkqVIv83Awk2jxdpXndw/8pXwsK32HW0LGOjUlf5ev6ETcsggY4GMOWkl+bij5wAt9LjqJ
bd9GCnM7FtY01hrvoJ8QMKIf7LxG/u5sXqTjnUbFdgkSRuSAbGEOXRJrYtO9kI6r/eDTZ73EW+KP
uJfPjEJQO2llx1fBzFzC9vcMAYBbQFZy2bpAJZ7CXBasQXWBBbV1XAAmCOsy7MZaruIPfSn8uWIp
vNK/2L0UFs3HV1mvSkUoFCvIJMEpdz1I8sSID2ua0Dab2BHPfZswi5twwS5wXAM7fM28k0G91QmF
H9svrZNj1Fe7OlTCTPQp8SPtj6pORw5zq77StXbKn+sFtMx0GYDtx5xwUh2SDXmqjxTWvhubIGz6
q8Qr/qiYai3IXDyGwQDqR6K9fWDzXGcV4k5PDyJyncAmT4bsmHHLEw2UGsZzk0uZZiZb+Yi1Rri2
XEAbxp/E2EglvqtESl5p7Ega6zgJ0hmWOx/6No3BWxwuzpmknxyFduhXeGH/ej8EmkLiAintuYRX
NG3Gclj0DubqOyXIUAQAYw9PrHSEAcuughHy7vxbLttvLYrRwPdOAySgE7xSA6vXVvNZ6Drl1RlR
yY1x1XldkO3KjcVUfT2hcdI3jTPUtIHHaATeOf4XaCw8xKJZ2W3Tu/BFMw8DMPaukBqfi5ta5H8Y
54sBv4uv8hbqn6ToriBx2a106jtCSa4HtdwcgGzlzc27MoyrHoSPT19G2FvpiKt9VkREDjZgvbYC
yl15Sym36HRCf2GeXzMRutk/UR/7xdNYwjdMcAFYW9bK276sovjVDMqN4MWT+FLZrW26llgFoTXk
wHYyctTo7i75y8VtPsWhaWHcCUZxXDANn5B8KhOJQgBTCAer8ikKepighuw4gF6Ep/A/xvibSGf9
MR+JIBGj5b2gWMOP6FxbQMaiMEBq9NBwYZfsVxtH3iTOjpjJiVIUKoX3RB0EZsttO1RKos0dxrfr
RQKv0Pil3F/zSdY277v93zXdbWZluepBvGdii8VvuwuGSth1q/mR25OOMTWBa0oJaCq3HZ4z8l5+
2BXld2Fvwhs2jXzgzejXrbm2hpsmuoqTAvC3nMnMc/WuQfM9O+WHefBFkxb1kWFZ/jY3XeWTePoc
vtoDFLMcdc0NTQqb30xRq82pHj3o5ekGqCI9t6s1VsVxSDgHCxTsJJ0vGFEyMaOfzHYz9Cqzjt5T
FJbDq+ECSnIfLjMZyhDMGNEDvw/+GdibWONIoSa9m0Ew0ySoMcVWz7opBbTYvjuyYJwiivWQVVoV
AuYi4KceGmRKIe2sNpcxlJkY6hOJNOhXYzOr//+0cFd7NEHEcnKh358T87orAykTpd+QtxPk1K6e
eNjWPd/C9pQCvLs0TuPsMpg3Zjohbysr1QDQOL29950INp+AYCxnpr2Qwcya7y9gdL6eVjweczqx
3iy7iNhCUXvHRc5DuQbxxfojbW0orMi9Otp0qxL3VCeaYWP294uD42CANrqiFYt23KYoSLuC/x9W
WPS/GyrQBWzqDzaJeXp1skehm37IUVhYgJRQgw3VTlygbpn6yusEl9AHRLeETgRXjqaI8swXuUfY
LsCLfyr8Xm7fU/DRvx9KEovJ/k1wwPFeLG1BVTD2zsblujkY2XLyv9GI+qU2z5T+wS5Wt6RPxxa5
SiRTqK67Bfg23FjZuQqcftfSrHuEvRJqXywozl+9SUwcp2gTAZwAwwY/8P9YvBnOzHlZb0T5vcva
XTE5u1WjY3oc3S5zHi02YZ/TR+vMVYUCg8bdKvXWOSerBHtBiYcIUeCDZT0TnQbAPDtgoTtXMl9O
BvPmo47D7ZtTdDiP+Yju74phE6QoJrNTBbJSEeXxcmO0xyiGvnZUxNaE+JesWC01+Byhrnynn10l
VP4uy4kbnT89/qm7Dp9S0RBopjbUlE168mwhP2d9QIFbqm8W2crqmE7sUchB3QIPbRIp+Hd/4tAW
udv0yI2xyfRz8iEcuxslWtJY5oLfRwSQE/9PqwCHZrafYBHpmdN9o06WixlyAmooLPuDaP3/x4D3
wRQ9ZtifCQZwxVgTbP+VWq3srpsOJthg6vic6tneF9sNw5opUuXLFBRWm1nxrqcdrCkAn3B8qTh0
LYclANqz666O3bGzv0WeW0lgrCTc24ezF1fCoQP0FfoebfivqOmPK+pY4jAWMHKEh5eDBPr/ZF8V
9q+MzWaBLvEO2TNw+UaTxW0/ZgXuSa2+7txhLi+rb64y6muZq9TImCJhWdZXbbWjopDgBk8OSs4d
a3rKqVo/H06yWTkKYBtFIgOifTP4xivc+KkK7KdV8ZjY36SQhRXCtGljpeIQesSgGQtVC3fKGmdt
Gz/aHFO8+VU6hTgywbpRHcIcLc+vtj0oBXE82izRhGvNNQMiOBMRGIiysgEsXYnQxCiWBdWZkXOy
CtVFpXkYODk5tgj7uqEoWZpCGdkAOhbVZL8wDajedioewbhkbHuzoFTyrG6vW+vCFFKwgghjtBRt
80ORjN0P+fWsUamrw3c/a8jdlvmXQ5jxEXDhwZPWpOV2RjHRP7XS+NwqyuhX9kkJHKdoPI49iyNr
6bhfFHWx22rHHzgZheiJ7uTaJFKUDpwdvJkw9NcF95ZpSWFDJJLfaGFBbGBhXfr77n/4/RijAhgF
Yj54LMkSylejCG7f4KDownkPZyO/b2NF6wFeTkQ+zWQoS6s2Y5Xu2FGRQQAyYQtCO/Xe6Zks8stY
yEKOEFL63d1lEebH76KK8Hm7QOlUv26V674oAebCfLv2Hm1UWEgX1NdhHFan1j+ixe3Q9NT827WN
IydPgBL3085x8+N4hyA2Zfq6A3FMsI3Gliey3S6h2a4yemW1J7RdKrSO6DFCa62DSpTGqyza51A7
46p/dvDp4fsxY6nrYavqlQ11slU3rb52xOPTvfGV2gbptwrPm3lMNa9P5vpczlp1ZgrsB9TV/tZM
dW2hf0O15HvDFiBcUI4iHfq4dDGpPxRBZRURsNriNzh00QOg1CAthkku+JNhAF7IJHq20cvR9B5N
Ek30mjLXN5C76wGGVrWvJ759FivZiMsV8rHPh021sJpcT41N770PS13SrUq7Lt1qU6/7o4ULW8qy
gJqqZNRtwIs+wus+j1pV5gJ0cHqS0SWwHJGa38FoKJXf/ikjU8fjB/54I3ZE67XUF997uGoqpG6T
qTqTam/aZ6aO9sVgso6AFRw8DdRI2DAL6crO09lCBSlpsnEeE3VcQAUsfjCd36rPmSCUl22xDa7f
l1+qiJa/hyEG3r3xFTVbHNPLx45aQhrIHdKvFRe1n7gd3un9tly6FTAoKJ/nhR2HmeCmXBk68l8R
BwVxeJR8KJtDf3sFYwBioX4PAfYq/zJ5WC2jji6KbrzT7XQzaQILxXtJ9b+EL/bWG09BdWd7f6+K
7kw2v6IeCQTnPnjdFQT/GzQt5jrBvvaXQmh89icgaYJkoPzzasLytOktZMwWtakg4azqGMnoMg26
W9fNfdr1CIFL6JwxFyeirhZfHX0rRj4eStvEDvqCB/GIvSiaPUT5/j9EzoJgQ6BftO3bfN0HNh6m
7Hk3tRAJ2oY3+ox6NGkaei9qeIy4yktj+WuJC/kgafG8khVVel2zwGV0xkfOgOy/zmkTkaPoB9xz
FgVsXT0A4Pa0eLCeack+xqFzI1hghvYS4rPW6hW/lmEWpCcxq0wS0CBXvCcOtXLbUozgPwm4Fb+v
toKGerq1kSCmXNRY0OCJ0chuygci6V7QvGPZlgVvMKt5FuVJrfp1Z7XknQhaUHh268pzJDzzr54P
4RtDyNulNnKy8gWSCAKAFfITM0FS0GnHDo2Lxybpc9UFBCd3NSSMAT5RvoNimLLMMgGkyq+eLJCn
YFOaiW3yloRuSfF4mHoevjIHqhEBhNpxph+vsyB1V+PlFy9zmMXNP6esttT1OgzaJ8jO3YiheGoQ
HFtV9sqvhmjnBWyLM044gSSqUwcYbY82PO7iWZH119RFzP+AlzRpfM8gnXdoGtvW1cX3+vPKIri7
HFbLGSQ21xZKfAX0c0L/H9Ocxrt8kkDhQSIf9tucFV2Doc4X5E+QtTPduEFC0xf+Id7I/vroDqC9
kbchAd+FSC4/lutGUrYVSP0noOOEDWmGmyE65jGnqFzXuDoGarpnByc9dwiieKUMQZr29EJbI3zj
X7s/ASeJSdR4PcmWw+p2g2veVoJOubagkPbS8OAxuXx8l0mGKlG9lZyiaY8gDlNO2E/uAWltdgGQ
1sU5F3hhYEOJBFeAvt3LWmz2j0c5fxbr/uLG02joUKCNfR/XKOKBs8TYl5uLPpFP13056yHlNXwe
rKcqFQkVeXjaeNzPzWNSVkMZ5cdWCCJWWBnj6XvKPYox8hn4Hp1N1jdgsh9fH0hiHKwoJY7EiAuf
ETkP0b/VBUacl6xLLi1maF3D3GxDFyMzK6/XNRr0t09fS7THznAHjqq8hpDqRZ0naZHTL0o7BoA5
5n8nBpCFd+8G4rD5zBNQpWyE3TLCYo2TPHmHjoIXL8Lez4JVrQ8lYt4yn9plITvumEozqF52YqN1
ITJxsY5lW5ZxhUdcea8E0247l4gL14rjoiACWbGGQINuSgfvfRirdVSU8Y1jxldXhU0/ljT1RUuu
X+1koFXPaLWKFX/VpLBIuQKyxr1yEyp78GJPLyVeYM3TmdQGvQ0ez7mocM4qZ+9NjprlDt6qk1yF
uEbmpenGpIL930gdV1VUlsNpEeknBwRn5uWm04fZvwW+uiklABGT3T340rcmMGVeLxl51mNkx223
271bltN9c5Od01PL68Psd3RxD3lY5o50tqjudv5ue77rY6v4OvY4Yz4SIzf8RPUtCMsPonRvw5el
Xa0tHadglKnSRaQ3W2Nu/driNffwpcMKLR+oDgRVvU0m/aib/ihYRPuvh6DqhObaHZzfp4pAGepV
CyB5guGBUMDCduwtrr/6h/8BhJd3H0mC4oJU1DpXuwTDdC0TCgqDTmn8v2N11kjRXgnq9z6H6hwt
+pqO1Eup7PPGUYRttN3C10ipz+jVU9AhfvPjqyeENXIOXClwL5/hSeGJCUF0UiQMGyJ4H2eXm6ui
1jd0ZMrgmXwJ30+odyKsZJ1Kgr2o3rEV/HeUolzjuTdxMxt3ZQOhUfBaLvy/idVm4zty7nqrL1Ef
QCaZzucYVxVSD8EPN8pRb/bC/PEfnfV6SLZ7Vll6j2+81osjzlZFVL5wKWeJKqwQY5h39uM6SAeV
smlVIq/12zY0eg8J4RFCKNmhDb37OtqPcHxjwYXJ/w0VYxvZEuK5DHYG7k2XtHrT0/HJQTm0Qpes
qdpQWBwQngpA783v377/lreMM1IfK496N7PJ2FaQhcerwUG4IyAtDqzLTWRtPcWLZhZHc4tNZhU9
HZXdsuYjdU00FSutl72pFCcDQMlcXjJ8Q5BHSn5Wbhmif1wcGK7N98/+2BS9I8PiPgBLH3drU84x
5W0PlTCeWYm63mEbqLqiigQfU5yZJjDvzkBUA1jk3h2XzuiAowjKynXig7KXo+RbSfhq045BNhg7
cD3kZA/oet5pyGsU0iclBwU5nFH4/2e0lUyh9jfIeJ9GY0dPF0ZoTZkndHrdSQ6O8GDA43wmPijF
Ug4TZTHf50UknBIpuHaHnFnLHm57FP3LMdSO18bMjVKn89lM7opVHyV/Nin3ErTN3bpIOa99DJQZ
QjEeMGVjHj+S4ct1d2Chbh/4meiFSqdWEPbU/oLJ31Q4Hu3ooVAJFJWz2X2HA1fwIGzUxtu+fsHj
04M86o1E5TRKpI4VtlVuXf0WIcVEuLxbJ3xiCcu79dkmSqdZX9ViBu1Kc8AgE7or0U6fxo/2G56K
SjEcpH0n/It7RyE3w35CJO7JULUQin5j3bpKN1sQhuUSZBf+f6pLL2D8w6A0+lDkXY2VVzPrsnb4
g3ycXs1uxC65KtDxRs1mFErWDvFHZu/Gay2VKBKYxKjT+RQOnOMTzWD35v52mE2RHBv5Dwt8PHjb
xuSlbipIa3i2vqkeGuImUgskSUyxebgEIWeMHHAqyH1XUpzVCuVLK373rtbDBKAIbaax/c/Y6Dse
TYaQDwFE73x3Lsj2c4O5FApICwcAvGY8Ee5T1Bu3aaswN7qtTV01siBaQs02rd3G1Sx5SPs99dpx
uKEFycwKzjRuHb5y2mM4z1zeKbGugy3cBn1Dd9dG4ZOvlcWicE4zrgQ4qCqzoPaBIqGPKt68v3zJ
Ouq2lC7y2w9XAoM4AowUKene1XHN2+nxmQbt2hXJCUP9ZsMeATAWvxo2IekRdMENvhL3p6BG0DWt
moRAWVxNl3DWJKP4dNL0C2tiaeuqUnrW0prraNYQ30hOfowiYejOTnqsqJQZabRdrDcVlVTGOQBa
0AB9+S+iwwMrDWHEGhO8ey7DjrNyid8RY1PmVDUFECUho9E1bC80pigK6yriIbJ3HPdwbxW4Sggx
gB9zVpyqplZAEhEb7ycopFDAO/guCSxd1OAz3F0cfISgY4PV6KascMMhYUwA1fm/LarC3MOdtrSq
xh3WmqZrQcmIdVZ5ZipwlNabkYC3LMPGhda8+ZgQ9bvkxkdkKQ1kTXsklENN0OFIV8zoXd9Buboc
jBML02Y0buHLFXKAsJXmQAyM9oaqCGocc+blLzLkIU+SfVyTjb8XhLruNpcDvU0gNiGxC4hKdsf7
lXjc0oa1Xk6kLgyNJ/qI1ezLCDuNrFYtfrEBX9h5GbSqxkXZAiwdGvTUdHeIT+1olhrxvzfEakBa
kGh3n82C6FQF1RUeChYBe9P65rgudukCcbQh8rJj7Wz35ez5XfSl/WlIbCojySuHekDMLEuteefn
gZmQekz1+xtDIkYAM757P0WWN9TJ6vQbmy11E6aIugWl2HJcdiSWrsuULPG/uFCkkYN6jvC84nCX
FThFOhXSZSf/HtY7+vAFgLAHB6MM6Qw6cupiZNBN8s3OSjPIFmQmc4uefeIm9D00m9tX2xdvXba2
5lYjDHO1e6TVQ+K52AU+7lniypvXfLijL4/jE1Mqh6SiM6U71+vQxWNqSL6CH8sg8cRb/B6pHq/M
0kBcO7s84IfFgPEk/Q2dW2+FUnpzPmT0acgzh6rcAAUPsIiFBFVzOkbvDKaKjXORyv6PIKnNH68G
1yV82vAiaEJq4og/p2YNhafFOSht08pGmbKvG5j94VCVJf3Al6MKe7WRkpbQPy2V/EYSNQWi3TDm
sh+VYxEGTB/70aneA0ozM8VBNBupftYCU6KOLM5q850bEt3osJXaPr5Pynb4kU0pQIPT10NCYGfk
9k/UvFrEWv2PHn4dI03sZ7nC4Oso57Pc9fNjeGQkb7RXVasl/t9r2jF/rg+MMCgk0EOlSHBVk7lH
okdHRJ1BC0dV7+4mLqYxoivaVA8meleNKI4XAViyJm8qricHkJcwFy/WNh1AbjyXR0uQL2frYYaj
yHNcccY0k6KhOFP6mFTMG7qvj+HVcct8RCTegqgCZ2bgi1+58L0jzuUGdsr8yxE600AmphUjFVxo
+bWeACFqKJof12v2fJSFD5NS3pI4FRzMxlTJ8j1Seuy9xkw1gjxkXhm3uD1g8/AN2+RswMg+7PX+
OcQqy/MQvcATyJiXddUF9PMd3AiNniphXy/Gz0Eo2jjmJpKy2qT899FhSP/NoD/i7zbf9AQ04ZWg
3kHgD5vGONVFOtxE497L4CF8fjuX8Yla5UmHPsIQEm3ridig6RqVipN/0loHFrM9EdwYMCLVFbOl
EgHHAW2uetfcm7JmF+/EbFTGwQgTTu1AVZvmdEJMCw/1PthDIjjpjvJWmdBV/QBn9LyxUT9mMh+i
FnDORw8Kk9rfhWy997qaaioPPYmjzjgTzqb6oj9GMhWbABJgDMk7WqiwOgZ390SbOMqdO00uCvVe
/SHB3d4Gh1KeKtiV6vxSISZFqAu5YMUj/6NTOH/g57j7WIRZxPpo9yg7lVyKSVHONMIgE3BW29qr
HJ0iHBUcWVjSNv9UHxVm4yTviXu5doER2bU2EBKXvu4yJdyOJ50JJ/CbpAeJusOM83AJPa99PDFk
S4Bhni0qcdvFiTXJphoSF2FSQO3QrsfEOZlvrRoy3NP6mTjBVwzFL4uCcLkww70ilOdHmJhvmLrK
vyDTQH4/y7yPJmUSuwCssB8M/wrgMDaWWXe5u3xCl0SlTV78Oba4Tnjs85ktWOAGb5EoLbnr8FAc
3g9n5L4m1qxlwz4NEFqrGyauGlg+66wXCIXUOWrjYMyO6tFz4l5gJHZYBSKeOgvnso9bvY0BDvUb
H+ORmAeLd0H5E3kGJ9Gxh3fCpnk8K2k8dejbHjYTNwwqFtOFm3VUWCQbKVXyKJRGGt8jGjF9Io59
DuPgc1hfYM1Dxoe6nXsq8r+pUNNCe7707QdU1vFumH/NVDoCWCm+5PFxKe4hASJNZ30++oC0sh/w
+wkEBji31XxRCactiNFH5yhG5g+TnBYc1rU/86gdkVd23rH3cDPTs9MHT6saU3AaZXCC4IojoAVb
s6uj4uQtmLuC5b145PNMGJXTxzCYAT468JOrUimQy9/SAzu+evqToKMziU8hDYpuHI2cFjAonwZu
EgSS9N7/wMb6MHJzO0EDoK6NjmE/lQXybjnFlqyPWYHJracS8vBs/hxEstjQOS8k0tI20ywTApiV
la5HASHelLbHJbs+EIrvWge9weEeqAhywZ+7mK3hYhbxar7M1FqS4EfW+FbfX++LL0MpBpgSPrVh
r6u373fy2s3YVIyes8T0TZABYpd6ifxiRKjXyN9iPV8Qx6kJL5oYulXXykmowEeG2Ct+xTy0jq4Y
mTT2xGMiv+hni5XiIgLbM3bIQ46gyw7XF+fW5Aq9UmI4FrPsFe0N9vpAcm+WOAP7ngPxGiJJkCGJ
xgJG8TFE8efrqdE9fv5ucRBfBPs7A7dBjam9VhK777kUvrs8cSR5RCOQeHcmc/eunb/Aji8XLiDE
FD0//3tqJ+SiejBQBzhCh8iw8NRglGORqgxtzQPkoPTmVUbjvzgIPAMk7eq122MWA1xHdlwt94HJ
fnoV1sa/8nfoGK/buoS8IMSQMxlRERq4WVMeLtdpeKTBuWi8OjZ5z94un0oTNAM4XDOKgGXWpH+f
WWhpQQKrZneeuWv62Vm4NJ0HVEIwOScrVT5yr1XNZcWZIiyFFOmXhNIV9OXykjsYLJwzG3fMfRAe
qfqTHuCWlHPLN39OzJBfAK8stmr7qZClRgIp8sMQKUgkQul40WjVojFFcm5AWROX1ms0CmcC0Y8m
vsX6sJ1J64A+pKaaagpbGn5ta5yfVV638qQdS3mtifYAfqGm9ZgTFno8jMWfmQO3u8KCK74TWJAV
sztDyyt3Fm5JR5AhFelvb26tw+JSaN/JjHv9irVxrGhRM7k0bUnxt3JpN5eFrKRQnlRl1Mni0EZ7
1W5tq1KEBSIMa/PlPF4NAqmdQLNM/LJqoFOcv8i1p6+tmQCpUDD4Xd+ZpYeuEZwN8P9m/zKV0MbT
NwEHF7ruUGIvQtWtQYq8gBVVdZIsqXdQaWxynAWu/eY3CyzRo6EXdWsPAfGFeKCUAqqTygVAvpKA
AEnW3l7SRCymiadcLWa4Hhj9oeFK9SrLW0QN55eSrJgs51yOuWP44NKFxUiDzCiKw2+YFhB5SaAu
zCSNukak8+GeoYTRH9+k4KSr+yzWjqR1TywqIErvwcCPdrZ4M1Jm8KxT4fvxAkJPNx1M6LKFqXe5
9P6wgrcF44YVjT0zU1fhslfq9YZoJdKfKu7KwtptusCp11CVgrt+Ux3pgVMm09T0x/hCYtI8/vQQ
KL14Y9qr6tOE7JH5NzR3VI3w8iU0jPQRYhj8pftPInd7Pi8oClnShx8EKPY2KHvuByHVqjnYehig
PAGscRfRLvFqQygKnqnIIOZF4Lsbhxxw2Y3zXRIv6dsw1WoNeEovKejppbcUdj8WPOIuMs8ca+ru
2XHIWDBvotMbx/94IqDY9/D9KAOpug20WKian18UZ9UlgR/Z1OQbukgCDkCxPvvf9MzadrN1joDL
7iAwmAggFuAoD9RtPl5NzkhtQShyPwEsCE76R8zpfBnsc9DVzoRS4VP7QY0aSmCg8WHmY53UJAVs
2vt4Zr4L03XPTPAM784zj0IOA4rXbxD9GVOmgRuLTpgyu4eQKWH69RrzeJRmvTIgPQAwfv2uHEn3
1XViu45rS/I9Y8LnqPho7IjiQMBsFOHqXVedyZvYqJMrqZzknL3snZKtzbAXuU3SkihJwC9q7v2T
7KIsputvyDKT2PHxVOCBnDOIkgYkC3hfB8Vg18pV4BbrRJsvQTz02mbVRNDcdPZl3n6opGlGrS5P
hBbU5tG/P5zmnnSr1pcYtqq1UHafkJmj/HwrZ+KwmXnCPtarF0Gh1YbyVKICJ2HpafNr6PNshTQ9
1CtsWgrgkkz/KDj7rbTWBS7hgkrDFTobJ+yNwC6tlvljlYpav61g789Jfqmf5bbqLdTWmFrd9VTE
KPcrSs5dHR2PYiWaEN4KI2Tw335ToMiuBTk/KLnOvag1ZUBFzU8DJsdL7KY4cYDzfmTcVkYIzdqZ
BWMb+pgC7Zw98sRisgV6EUuoN5nIj9GFBsB6/ro43LEpW0YgC1z9gZZ9MJbZzeqvXotw2qD87DQZ
a6dG9r8s2LuOlKX4lKIPuadd9g0l72H1Ko9OrGnUfnsDk1A7VIlyz6jl7O3TRKFyGATlU7R6GnDG
QwybBZ9WdcgMnt425y38EYBV95lGfz2MyjgtVOFbymNB+nGA1X7UegywLYPNt3bUZyspDdstGV1V
286ohC0r1PGbKmLBpl3s0QQ/Z97WFpz9/CPgBP6upNI3LMH4aSUmUGDS8mO6JCCmrZ8vKHdE2Btg
kn6FwNebrCrgRq9A2mkPM708JsHTOD8s244QfUcFdahmSVinoE7tODfwm7pPLkaaiUOvkmMGsqSF
tiLDz/7pPR7Smta/oYUuaBXIVKYsRioIICgNDm5IlyfQPeM0MgUjQ3gJUo3pd2vMs8DeInmIrr11
Ncijd7+Ly9sGtJcgtfFCe6x2qCeFVh//gbfqtrjXcyeOaSPrXpsXPUj/FTPjA/tcJvcqYTbENZj0
AKCfhNHx18/Yb0p7FjCVuAsAwW7CtuadNHknE2i9yTuA0Jn90VoZeephts0DWSmRv4UFq7iV+988
lyNAYOpAEThigiG+b5r66/8CjboNmlr93J1BygwNMdBLdJK4hlCJNmyxW9cpe2ZoXIV93BrtFRp+
e73sDz1Y80BiNmciQWHx03R9n/5LiOsqvmpOGso2DfFhtgis4KkhYYol31QEPoBd4dO/pcfDxh41
QXdlteiwcGSbMaT0SIxC1uqJfufYZfWJOstbx1swRKcojm9u7FF91aWUyLyJCJJ0EFAmBIrMWqN9
YmX0aEVB8hBuDNIXjPhaBETNwsToyQJxaBODdDU9fI6hBOZ06SlNuGPi869qbD7KcCGavQY9bVnM
W8TuP9hHFzzcmMiygB3n+Gjkn/vJCLzc1wQH3xI6Wt5Wz4H/8rIntsYlJJ5G4CLEfrz4OXJV14Pb
LMCWKJxPllmeb58KTtw4ydJqHh9W5Acb9YYvrManEHaGSia6bac/3S4CUQyVefHWhDPr/6vbYVRw
XnP85BGYU/WwPbSrq4JblGMckE5LGGU2Y/LcvCGf/Ul+59kLwS2ueuhNScOUGYOHGA4DZGAwIjMJ
XaPtcMbCcfJzz2XRp4HEZiNkpW+d96g9Lir8vDuIb502ZRLMZY8WhZtxQ2cw9Ph1tfo08/KbaQlu
8gchZhArdw7nfpLVohkyKP5Oza69Ay87WLaQEkcfGQEFe12PSDQePrXROFsluK0T4qb30NlnnW1/
Owc/6hxt/dpFGrPU3pplLiycZ181n4sKW43lshPMBplyTHj01uAyrWJZVPMYPefODdmrPjowJ/NP
+BUZ3zOPdF82LB22CtbVbICJ81sXZbMZCMDN2gLqmAKDPUS5lIm0aPSoDaJUXt2OWlYJXq8B/feH
sd9PKjCSlxmM9KyIhroAw9zDQWy45RkCjwNB6ypNqMffe87cp+iHgbwGv3HwQL4uEC08klP6K+nc
azEWtlX/AYjOrwe5c4/8GHg6J20FA0IPMyWZQjhGsAt6ywP+W9bSpz72y7+zfoVUlwXWGHdH608w
y+h4c+9EiA+9kTNbOGRJypNDe7MgNwjJY/y6I0ABRHEd80KTLJZoMGNkVSJYYvmTnok81KdUHi5P
dogHbfCAHdRUYMr2bLt+DLiplzVJgL+RLrgQhMNNaele+jy52NGjMmpDhWz9QjG1UTLK70nqAwu7
gYuki36VhofMKqs/RGCGMo9Wtwk1rdG7gxoW4KZH6sOQOMOZ6T5DFLKmIlLHVv6ML4uc0ojjCxma
uZdGDRUDpzSJt7a+XXLIVQ2IxvbyI30kdvyzjEdBUKVsg+kC2zs9dL/ndjSkYTjMoZvV7m3n1CMy
VUNmw0SHHfqWS7wKyrQ+avChYP8v0tMAjY/QpzXcW6c5u6yvjvVgNEOhwkvW0iWfIMEoFR0KdY28
B9GRwFJximgoqht/wXKRX+i0XfMml5ZbeqdPj6hJ6gIofIuZB5UcNm7pc/Usoi2Xel/v5N0RVOSF
tvqIbYc0b5gAn9xuZ1T2fMRfgF+lRIfzUV1goOds6B9ScHjk2DIz5tyOzr9Fn3UQVdts0UC3/b06
/iEHSX6tL/2fNYrNTluHGPFSAWNelBFNDixc6gmNeqfE7wu4tJnMkWZopTy+SDSVUgy81cLsp2ij
cv51iDtc4MHo4pTzlAsn+5BucrPRW3KG8KQSZbI+GCjvnw5MbzgjbGzQButEHzcckfGx528Ifmfa
16b4RCha4W7ij++zUiRRdNFaMhrxfZJVjL57jaKCJFUBuU+0Q0gSaDLGZpafrHhuewETymJoVyaJ
/IN1rw7984WI5h7b2boHPsDYX1SXm54TeRABLsc7OZyGouY1L0wqNhFh30t20gy/9BdQ1tNuzmVO
4f9ZOKZp3hk01drLiT5vJPxDScSSb/UuOKiv1W4ajRIW+ziwHJXpOieYl39gvdUx+btZU78Ef1dW
h2PLWsjvDMbO/ZBhst3g/BIuP90IP/LxtUIGX3EIjiI8z/CIpwFJHI2AGQZQdu4DTFDq2TZvBk/Z
dIp0Gqvg0a25uJRvsoWdGj2j8/bcQleayaqtCbu57zS13ouns3S27Z4HS+22i5+km5SaQPAb0Nwz
UzS0gChzKaTyvZ/NDEWxFNCckR4NSaPrubOOkE9qC4GWizyZ9T+oMsMBrp6P9u3pG0CYXq+2Raml
PYlCJTk4zZNMdyRyg3wzwXwyn1itIyEaewrVdqDciJxeJMGegY7q3wyQXIfX8vSy0g98wiyynt01
LgArRnp4Y1fH9avE4AxlrAB3lDSdbLucEI8+w8mud87EibnSALwK6KDzStKdeiafoRtRF5G3ifNF
PGaVKw3TZOz7Cd1KfR3+sCPC11DCnT8IE5vk8+tqbklU3q3C5zSyOMB/k60kDyNffp3DGtK5gd+E
o5FC7GwCh6iKdLndSgt6Do9Vzd2UzrsKvTTg3ZH5hSBmyoGDf3SCZvweSOGWZpHKob/ETYkbPbNl
tJh+mCMb1+Vw6Vd3Sm88DDoDuyURfZIy33Yu2b3yNuTd+ZEk8bfhLSYAPethJl1rXGLM0saMF6wI
XbprHl6I+SHtWWEVtJIAFccpwK7wFvvOSR8sVBn8eDaUmNAsUX8aJPy7RBryYV1151W0MR5X0ioW
sEBpOggRWW+0WAsRnnK+oyMUveLiDEF44VhX/264z74I/jOkwSTqjPAACGedhjOGTJCWUmHB7I/9
SOQg45cbUfC32Uuv9+ySFq/OBd0HE3v0tJKc8eFnvRKhV5XAePiRo00Md+nTE5X+tIuTlHSvamlX
miYXHkC7E2kEalhKmTb/+MbStJWfDKX0wLbtbC3Zp7tDRHxudQqb+khv4qDF6YbGyf17GtILVO2z
7/jFLMHnGu9Y61VXvy/SPjQToKnbIsNUoYEV29vV9fVLL0Lw0fb406Hx176fCDWWxZfZwGBvU//x
FjHhhaBX3bUoha5WVffsthnbKRhTTnSdBRz2JiFc+bFmrrYRcekgSHvHpHmCg+8mvcbGyfpRfLEe
CC6dNjQiDitbQOu93fouwoF65r+wdpNxSJYLHp5SuaSafhr5zz9p+wkDTDpus6AF0aO8nLAEn8Xb
JgvtoYh5lcMzYYoDDdT2/abRp8RGmvhRB7OBJ5aEHKIKOO2SmTdpkqbFBRckDttLSEm1FUXHLKqo
TK/1ojQCOJt+GeGSJA+Pl5drW1VxC2ijgnptgbjtZMSvibFPYO1qRXIqJpxzSI9FLWMNBj0rQTyY
5e1FabsVsiPW/7GDor1bCeALiQAQznngPvGrYnvCruYDv8sIdGtl4T70uBYdVdR9g+JnJm4WSOzb
3v64HZJ3oitbEAM9xJ7ge5OXvi55g5cMOlfP5zCU9qdd74TfqQH0UEul1id/09vyno9OOMbxAsYW
46wqvow8d4hErP54dcbnyEV5lrMXTL3k3MhdKhGJXc1P0Q2CNmJaclalOVxJOBuO+zDAyXalxUkw
3h0yMFhJ7K/xY1g+UxB7KwK5V8czY4e0dGgZRWVEf4bbOc/XtTl0Ivw9TZHIYYds8+Y1kafNP9i8
Pgt5XqkmGJpY/LyaYnQ4PaNZkzz5dhoLWyG8FCSx3x7nIomgDDYxyr0FiOU5BLa99gGYAL60FMMx
xqzVLx42+B2aLAI9Km0xXAvz28pi2A2KYhsJTJCrwO30T0edLl7iQ9C3ggeRUnfRnK8WE7tMjmbA
yvCfUnN6+I/y/WAvLn9vAPsIJfAW5MjNeyHXG+Rsfh2/7t7sWpsFUob9SM75qd0wL57lm/AEBL4X
3AuMEuvPSasAaYur+PqtCXxWDj5QE5HIkVvoPe3SPf8Fv2BO9nAjLmb4Gwndb0BQ6XK3voy2N0c7
esiatXRIiGmDEWYBULnEK2lxXUTDEjUOwpWhXmz9WaCBPuaA5XmL8M1UjX361TCtg/LBNyLT4iGS
SxSdr+GgjdnyIj45fKEH0icN7b466wht1oKT0e+oHkvuE8NyvR30bfvXWSVMmWcokMyLv88slbdW
Hp8Wny+6Ba6C/RH3SCyySacNLOXv9lLxt0jse6V1SwELMSkw64wHi5OffgOWi3aGL+satbKFmQmN
vQCUI9mBhHxNlY3NSHq95EmZok1SiXo+8jB2LloiYraCbg+zKx8rmql1UYCzB3tsOVm2PRaVXLhb
FqN5M0Nb5mMkDA75eLJrEIlNQoeXxhDppzGbVvGbPvrBq4Ki4nWCl8Nlau1xQ2qau2MoxLSc80r6
BOl60FBpqwc56+A+QVtuhW9BLhahGHwOByfuwi91JhakaoZSEBCxHsBzw0fNSwvpo18Z1bpLuJmi
y9YVnEXNqG6NmmxFZSa8EwK2AbFUtNrGEhueRsWSImWFBqchK91uV+FOMZmAnyAyPXqU6TgtmL5M
zcbmfDoWy8PdEbCKhJTD934mjhRGFsX/uBExcjXWtlc8lWhC2fmfLVbzbgV6etn2inu82U8IkSdG
1x/uZVqTNqCWZY7+brgIkY0S5XaQA5+MV3c76TIGRFcbUzHwwRALzIFDgsIXnh21kCwT7wRw76DF
10UVuWGh5BLyiLVKD9vS6cQEOIw8TCG8RKAg7zF6iVPby8b7yTUHVKuglX6sTmAEMueBqqan63SX
+BeNC2Jb5V19dPc/1TdL8cePvULvpXq/S5OMuEDUSnt5+2n+8KyVBBxgJC9AT9Lfe1vM7TKMr1Ga
zqQbzeq7hRGsWTjyDaF5+isGdBDMtJvBQsmAsZUEBn5/Dn7tzsH8qwhKcRdGOymgyIPL0qHkTFXM
RDPGoVQqpXHXa0VZulACSWltkUv0i7tpqjrN9Gjkca41atkkaGgLflJNAvUXf7tK87ERlyrmY4v1
eFcJE5Tns0e7fz1uxJy0CsRgAMnRKGxFlvYYaGDelqECWwA3f1dUxvI1AECUKxuu9sae0sYURFaA
MCt1IyUWOXb46WFTiUbXXeU+xjchAcBCAgC1DITGAvYbwxrO39o6iAJsegsgb6bOQGzWS4b1TP8J
CmicCGzOAdykaNo43Fnr09uGkF4tdtnuaG8HGB8sO5qOb/saor18/q4OjeMnPMHCxVayBE60Rilu
s9aZ9TLW9F9R7LOJeeJALv+/efmlvQ4YKHc7CF5RkYMYIzqnthQxVPToTsBaHAUj6AP9T/oVEPP6
okMA8Deoqkm1N15kb1nlCVQYvELYsBN9m9m8lTwYTG00n33cuwXZRR0gpl8Etwru/jbY2l0wkGPf
eq3ToEhO8NYWgs7TcBu5ju5/PvEqbouNgRYG2QIne8oL6Hak9f2yKDo/VS9ILX8yFHRglp4A2qZm
ZAY3o4J9jpGKKvj85/2LMRHNNHmeJIjkv95J5X8l2dvLihxCK2ZftZa55a7htOUgcwRp5dGFXzwF
p1phQB7PpCpuxp62mEBtUFid9ug9tYu5/UoBu7yBZGqU4XoBmzHfL1bzC5/GjF40a/adqwJR3OHE
Nc0TTorViGEdnsg7qTza9k1qpFvdS5Wh1onyXCb+ke4y/Vv85RJTeXLi8C3GwyeUwwhQMbba5zIB
w148uqFThgTUI3NvzTxKEWWm7s2KPApvbCA/v2+xoow6fbkhY+xljsmyC+NOYRAAC24dOhHqlefS
2Ah0GiLDA8UNMnJ72ow7vshNWp89ZGgB+qlP1Mdy+pUbralSkX2/Cf5AXeezT/nQsL9+/pIj+ZUr
//yqkMQb8Fp04kk1oHK8H6Pv833EhSltsW/MgNJpYizkPvuT+cRF3TIjg6oAQpaWzI23eF55RoXS
6AAahVfXNEHxL/vtEH6vy6AWyKQHQcqGnVHSYMaTF3jBoCZSZCk1dG6puQGWC1kvgn5vU94aWgdB
tufV9cN9YrBKKmXDc+3THSmxuvDYD8qw7Nb/zks2qySeyLYbnSftDdNiXMSpxzFxnB/EdGujKnfG
CnKOgcXb4g9Ai32VJrGmFhyZB53YvH9wkhwWcqWR+AeiKqSPMy5DSEzthm8vmAd7LzzqjbjeBQ0B
7aM8HeZ8A2uL9l/lL3fkVGsDUBJnoMCpUpfCwER/CAkDakWc3uXVXWJzeZyIGMa4f1OdWubdSHqW
JYr7FYZzmHT5LSAbOJ0BUkktJR8YvF9Dxs0RiToYVUtk98h9zFQiVk9Tlo+F8Ud55awgNxQMyCRI
EojdBCPyrS/OZKb+Ij92BGsgZsEiPcNUgW94rDiipaJ8eD9s6zMpc65JJSlKO858cBFeexP6RY2U
JKDrwx1FZz96Ie+u74V/8/tr3RWFvTkQnL9rnhuB3TV443dyzcKQszV/BGTdcFof/8uItrzmglYF
uJnGm5gWF7OxEZ+rOtc5ceM7Jo8IdKy8jG4bkXZ5/GdGkhDezDR6mKm5tJF8LtvaCtUFsjRDWhFb
4e5nBSNobUmH2V0wrpyJYTWpUpN98JBx3z9tQuyCDzIAy9o3KGht4uicSoGMB1dLap3PsamLqH/p
pCj/TJ55YbeqwymV0nKWha2iS8uwQGlvhBHWURT7UIIADMN6F0+fhoStLUEsTWc6pXIobhcA30iB
e8k4jjmzpGSkGnBdDjQ8lx2f9HdVZWKPIxuDy5FosdlW51/UP+IrEq4hbPKQumI7EbWDNbC0YGsL
u0nEPUjpktkfXHl07/Y0vpKJE/+0bWXDUnzMxxakcAlp4Qlxjdd4xhaiVP1gMk59ni/+W6uWU4z7
2WjNJwZktGyK3E7413IIibfBd00g91ku9vZNftuqGxXC1ixFmz3HTz7a8aaqBf+DZfcKZ3ItTnpA
aJd1/r8xixyj7DXLCvL84vOi4foOdEUfd+BD5yzvoZ4ZrRv6dS8FCopNbzlQxeyTG7cHQaFo48ol
w0ym4MXy4ZxBkd2g+9iO/A2TZY+pqJN8bOmpQDbKAylNDS9SpSI+hs5CP5HBVGzRONdw5SjS+zWp
rq6mqDZbd42zjK5iWHnHRqmR+/ThY3AXzXYWsiUZK1MD5455iRszzFn/I+uoAK8yTsgh5cwcMJzZ
WpiVwPGjipSStXavS6ujIAmDZHCt+ryx11OggdB8SsJrijzx6KLOHVbLIjLxm+qBc6nBIvrq/0UX
B/I+zwc7o3rHVBD3eF1web44LP0HGj7cX60Y4ZDVyiLlCY1f7sXGEkiesC4wmzwCpfrYlZLxqkbo
jBwux/xOtg0YwR+B2QFEmB7oieku9aAkTdtE1+wskwmsYRRD57coPzldd/84JmNH+qMQs3xGbYg+
VFmQj9D2qRg+Sma7HHJDIIMK0FafyBqFArKTbUOcAxUbXYyqHYGCJwC2l+TpMGqCj8voQYMsqgm6
xdap7R16HBhlUQlqN1tSjaEeYe9q3NhQOjxNdDo+NVksBPSggjJ4ZmodYN95rQoHK7dRtRnKnlSR
4/JLzt9fN32G8RnacS72rvliNkB4iirMrb2r7OZVkYToa+b4Tw8cR0lYdVEzN3Q/WqYE9sFmgVQG
GeW0kLKMTWoGScKlEERaXupg7fO5ktCPrbZqh6NhJ7HmxQT0G3x3p7imsmPz6zAzN0QDhjHneI/3
EXRXbGcxFp1Qw1Bex+DOmpLuYbVEzKrdXpYkd1WP3iY7xDQkkIof43bx2/WbWP4vdYfrTwEmeigS
pJtGawVDbvObqfj7j1UOnPcKHju35oRNjhNgjNZ7a48iNb0kIDPyLC9NwYHHhfHroTS2m2MlK0w+
DOzj1JWWKIuuQH8Og3+bGMBPHgJJIXKN3GeTNShd9Gh5v1Y5EX/lvcLnK9wjMq1mtje3YnFH/iCT
y6umnw1zR4GEijkygzBYhO+OXW3uDea3n6zuMvNfjrg3sKIBJhrX2L5HrIjoS5oAy0sr+D5N851I
fth9mGbr44zLSzy8YbWF+WvNwLlzWh0q7lKdeNzAXLLZ7YTcD3I9viuxTbviFhTlcLz7zh1uIv/0
sWPcbrK342ChScOeOEXXdd99kQL+Ah4rmk4uyyC48u4bFonWKhTFbIlh6Nzoemn9vWbqoc4pX6FW
CEDNYd3ozEeQg5vwH/VDWiBRpK+E9xxTlw9joy2v3rfdoa8Lu8u43+zsrNTOtYKo6iLr5MTtXQrT
ysbDv64kVZ9S8Dgo716ARlJ/rGHsVZimBFvONUjPeZAV8fvOLb6kbJuNa3/3FXO9bZXfuMP1KkID
+aBRLypa20K+RQuxFfUN4GrOZza1WdWDyCFaFYA8r0uvvn/0HMy82geqlNajjlXTDt1lqBvE53jJ
uzhiGklHxsrWhJvt67Oi1nJ+sRMaZD+YDCMTi3Nfuv2R96YDWl7WFGlZSjmpvjqJSVLHoUZm1vC/
vZPfAbY3Ix9RawijAWNDw9x9QLRUEb3gpcCL+mD9Uv4NPIza5cWVzors42K14KY5xznVvY2nK/rw
3CaiC+1FyEkoOzEQoC9iE3IyYAEoqFEj0iQ9Y4py2VJtzA89ABYtHXFyFuXoFSXG+TziSEiALJCd
lLJ8FYQSqIuBfxYKUPmgJb7GvvCzb+W6YktuLBVKX+6D71/QLm+dRE4D54N/uyOR2zJMKTvUWxo1
QpaAl0jFfOVMXZBE0KZQTWB3H6oyj9jRtu1rjV+8aRFsR40bt6Zxe8ibSkZ1ajB48XR/a0DPbARz
3M+J1KeHRgqcAlSnu+APzYH0SNfLbKi3fl/h5a2EjFQt2GU2/AEqUCtZ3jbxIMojNGNF/8AbF4hd
+WfLprdz6Sm1sNrqcDPQ/P/hPm3IC2KM7brZrGgKWR4Ytt31cvn7ID9phrxGmx2C/NTxILeU4MNn
dTnrBlTAO5qI+8R24ObY/ivPKHsfBCYztvoAu9/S/YYM2J4k6eHAFgo8gv9ypo+YL96EWARZD+ZW
B2d+OYFoXmzebmGhxSI5zcN6VNPYv7R2dmjAHLAFYoslDWVushhp0vHyuE4i85SjkR7IqzkmBgLc
UpHF2j3yo30ImktekCRHasmNcFx/FdmQo8DNKaHoyemOwgY6B6PmqSvoElzKvHCfSNt/zt0u6sbw
Nt9xkNVC0Do++vfDVoy0Wqx4XykZW63v4Wnhsk0nK9U3DzYXpIPy1yMPj5A+6FTtZ5kSj2JFn0f4
qvZhmMZaV8/iV/fgkqsKYdsrmnmzTZdaNCHCVRzxy1/zvaxb7HrTuG9Sup5r1/CCi1PJYoHJ7dsW
j3iJ6nal36++SfdbGXzI3w/MR7OjaErGt1KIZf239gLRDlEHVP1mp4NOkvojf+oR4NyOOYq8coGJ
zlJXSqOkoJzvpi/mOv2quC/DJqNZTm78X8A1pLqjW8lAhsQ8CAh8c4l3rtXz6Fb8u8MkBjIWDN4L
/w1CG0P8diuxkUCJ57BJCZdcw+1AuVBAo2lQLmDFtPdde4Evnd0js3Aqp9Hj6tMznc+mf8LHjYNd
3G/Xb3XNcFYbq4DASMdfUqy6l9Fdgn17ZqlVIbsy0xjr7hYZz7rj2nmqKtb6UnxnNX9jB6A6yJPv
OaeQGVGUb68SxMMW0gSXfmwusU+9qYDqWKw9rDROsL8cjq3RZxNMgOej15Grbt+wWoGN5Gb3PKtC
g2IdPLAKv4kzln6HHk25Tga2SN9Rbhg1qs7v0gVjWvYJjTt2/JepJEudp4Moy1H4tP7GhJPVJkgE
5bIgj5UqDzKiiqkF5hBDpOixV7atSC5MZ9Wf68i3PXq0rcuzUSEHHVn/ZXP4vmfZbQ1bZIYlkhSM
CjYPKyilUm0TTGvLAfQD1Gvxcwvoj6wwjkcpFI/pAFOBSfuXgidjb0rQq5ANrBy0Yzxt6E2hG5zW
xwa5Dr0saTaI1fubkbVFe3wGV/pVaTuzUZ4jnAHJigbVWXFq58e19tBm++xdWTK/QgtaOAXfNiGx
TqhzKrzfdYMmpERo+dN4XdwzwjHusnYbNT/OOLHo7XPYq9eJLSieVxeIzn9zDe7tyWxnOpJlB8Ha
MxQQ/faS8WOYSYb/XaCa9aikt6dlCpV9s6CjWYm5kMlWXljluxl/kaLfTnwY6UvqZyF/6IaciN26
pOJzT7pM0JFt9d5FPIHzU+vHTt9dsfYvFaPl3pjt5p4ucA7gjBCi5NixP0uQFEqyxAC/EYGY/+3g
94Q50auHlID+8/ZcZ6SQXPrtYtafCRQtVSZWWhrIuL8H3pwBaWtmdHkJN4yb5mWzlKQI+ygcUWST
RWyutYSWtv0Ox6RRq3tZLhrZFHF5DiiJIbW6TgpLuu8cm4Y4TULE1p3w1pTbFoB9QagXGcbFUSMm
TqqUqTvBMorZFVd9exqY8wBOW4k4E0ri4+VSesTKnV7gSO8aXZrw7R+5waI2jhd25X7ojnIl/FuF
yB5pgaRuqiNzLjb9pjUXcXBUGHaNZQTGfGffwn4mQjhGVVF7nNuCXIbOaUEytjdZklz4469hx35r
DAXSvbyjHWlKCR++nDOl78OblYz4L+SOJ37ASvYJGxm+kD5Wu+puCSBabluuYJI/Tl3Niaf3qgOb
O2sNIdG6Mk4Ti942JsBYaUEjm6gUX5C58dXQ88Z7RnrNFswrKeFeX1lFI5+dqouEY40mQVpy+XV1
yvgxJK5raSaZ2djpWvP+oXP3ASBikwTit/whnlWC9wgQ+ruJ4tyy4yCpYbN28ngE3HKgYXRoj3Uv
H1K510btwjPgLPlNRDMaMHwLxnFWwdNEtEwiXemGCI4HfcxHZ7XFOLUjFmAsf1tF5Gbdh6Wu6Z1m
SvNHd1VEVAekJH2JBN4M7QIy+7/upEkXjZYrpD1FyAbVliuZNL5Ycqwm1X+FHTjyK/kGEAnvRe9u
xFugHXKDhk9WbLpyFpBNS9i9C+QNI6ievEeMgf0QGaLeYrGQffi4wiFxSPidACoWhH2RStiOohYx
176PabusmVdaD+WXvvIG8IRQaK8YOwHT+uFVuMRQTh81UmF2b4NQdgbuOeoTdKRVnlszzYove8tf
cKih+iKvKwRsxnIqWkBV8FI9h3iEaH/9hGkqN0nnZ/Z7e0mzTRudJUaaL9OEyP5b6cnYdJg/Cf35
6o/h5mHSe2yRPwZGJ2YhGuZMFnDd+NrrmJdsPKnsjno9+lTvRdbeHw1wLUsKgMrvrJj4y6O4Dlcj
YogNwUmref/HkZHYnE/D97UZmpkl81yMW2s/C9OjKnRgtuPSKzyPprdtgPF06OyTzcggu+KCEhKT
Yux2dJlZXT9W/D0GgiDQcKs7rH36sKC/yrkDFkL0IONrm3/qoWN5Fxjq0gevq0KTjjGHgq77zfio
7epCv+EG66jmeOpzKO2UUAF39IbmS9jard2hdbmumTnz9HAs83jm46EFMOcuTxuZzMFCD0JjiR70
2hXEmeTQ4WX3SFOT2R06MFwVHl1XNGvISiJYJPMu2VKOTVU1tX5A1W6aQnaJdSC7rP/lEcDLHagF
aZM7IE1VSaFFWwupZlso0+8ysZ7FLKiHEsfnkLoN04neqOq7mJOpdTJJXPkyD0sbeWVrVLpHEnH8
0FomeNJDzb/bQjpgBDlTJtMJVIuOkbm514UZp3X9TAK0p+eR76aj++nFrH/VdbaR+AcM3rkPtPjN
cfG1ZuJlS9RczspHgNDQqn0+TQFC9nlr6STC9ybefEhH1JcsxihWIApKY3gwHpa5a/Hq4FB6qdv9
M6oCPLurllonmbpstujc3jY/RaSOtDGsHhZRmHX/l5rSO6SAjEY3K2GJOXPCpwu74v00ftpweugY
ALXDYy22tEqVDt+PSfG+uaI4CQeLZyvwUzWXo+9pgb85cy+aGAq1PrXb9yYVdfbrMWwQ5QYefYhF
VFC0jfg5IepXI+1EDfcjj/COYORC08zN8OvyMTMFNm/0PYD19izUz12EdbGTxXFkKc+2b6uzwrt4
51g5VCvtNgCs7CnzEp6tHyoL9Ynl+fa+3C7g0Jewi7x7Hj2X9SxXh/MwXPIC0+MnTsumYJj02kh/
GJWLfrfSfzbZ0qjtCD1OZ7XL69iQSZwqS7AV3SUZNTYnPf7s7yS3r1WQfZSRGmt2LSeJ4lNJhR+8
q/YcdvvXuDpzbmS93PdnRGoV7B+sfrAX/HrRXGKkxMiEMLyspTNlit79TlV30K6aFX4kmLRHom7d
MzT0kWq6577pTp2ArVSZ7J9NLOPLKrKN8yyYk6PE+2yrfo2Ayq1LdSGukb0BCNjbODt61DNMU6gO
96rnUqKR7kIFbHACxGTggxezLwFLVE+laTyf0qo/MWcwtszDb7wq1H3yifMX7vWxld6jV7eNEtgi
DGKD5LSf6ejW3t/BoorIOKieOIdKZ8jAupyZCh+Xwme59ewZcYd/A+o2WJB5lIcMBqIoMTAcJmEr
zyPL/cxMHtXXCGJJ8WdQW1HQ6ySvSAXgiMM748rY0w/uIvKxdaJYxP1rcLNfv8f8MA9dx8GfowbG
cyEdfq/fjJyBHqFVQq9nu5wOVB3TvOJOsG48MjS6y5s/da3K5YHuL5Rhogljkg1UVxRObMVt3jla
NIneAExQYw5BXH6b8Z9Wcwk4V6A6IUCIPTfKIfdKexotDRM0Dmuhy53rDTi+PXn8HjRP4VSW/FT3
TLbWPIgCNkLmLohGc8UHK9xhdGZ1yn7Ca7lt2oTDyf6hSBJr0tUWBg4DctKCH8u6v3w6FBhE93C7
2NDphWxlTUnnvgYjiPKcAjAQ9Y8CvTz0LvHaezvOnu5viKrXCFmTDmrHtjH67DT/VHr0kvOpdzyC
hDTnFJHEWNEtv38ZHdptqTnoOoSFePVs3egadE1D0t5AZOW8cILDWMjQBP5+VselEVOtWlAuGQw7
OkwWc6thy96/1T1uShTo+x9N/xf7rTBnz1LJOm3dMYOzZlwkFIJJQd/GPDeX3xsCBDb8ZZ4W1k7N
sTlHtFeN7CKgKiQ54tn3U8hVu8qvBk8YhHRNIpX8y0jAwk6yhu8KvBPhJO0VTJqZU07MPDszUuUP
kH7dtcbQCi3pemWMhKxsaLLNsjbhuVD1pmDZSS1WTE5/WKh4GbrE9Wt1UDtpwnC3FTp3ibtwCwtw
dpHSsnOFC+03PZC26B3Acp0xUZLq20rxp4oB4upmLAZjjSdLKOVEY3Id7qHK7hsegpDt0uHfoivf
4qDeSkWtUMJT1XdFnvIMQVb5ziwuRLwLEUS2rTIrvSA0o70jAt7cl3mg3mLNoWdcKw7wdRxiIjG7
zUx9zhPjrNbOybQGZ3jjsBbGBjM+OOIS6PpM6YHwJ2AYfkjRh22P7Bu5X+FqdmZAAwNOhiEkkK0P
EzsGnykXmkriIVkrIzWKHF3mfyNWBjB60Nqi7WnTOwPVoZBlKGyD7wVUOEKDAeiRTQyaq9cq4wka
8oGeXC0q7eRYsv6XZgeA5C6Rh9iXXEW8u7qMS09r9K/VZujDtbd/ewfTfIEgnGLtZUCJjmjkxn14
vspmixGuKxGXLmAsuUTbgtjl6BK7uqgUBI5jQIJdnh5KmjpkF5rTPb6mwKRTuBC87HpJmDuXtNcb
GlvhsTYHzRJabY9/JxarxbkjUDRNgID+phxCB1BIpg0oQyANplr2fSxGOyw4MUad+zEAZzq7ZEa8
IKcz+lGFCalrYriqgC/e/3YIvZVdVWb8RGqyHyxQiTsL0fnEDCH2jCRUQPY8beqOQBqHMrPc+Xaw
tOfY9AKs3gJEqdKfo7Rm2msOmXt2KMQBS81c01RnsYvvjEDsdMsH+mbr+73XXLvqGb7TyNXe1eZR
cRiXw05LbLLDOt+TCYPDGgdXNgyz7BL6urIXU0XRr/zZ/AgkYE93gt/d+2WxHPRPw5dhKDSaO3K+
PeLEn2TN1EzgKcRNig4TaGWEUndWAg3g2z3glFcpYHr6mMV8mjg7BEhMiHGbHLL1numN/0FHReWx
k9TnpFotTTwis28Jhc6jfNj4XTnR19GsBCmjDAj2fQ3gkYqMfyIOePtJYp9j/DgwMDoLXTbmxV9Y
i093U/nLGmnDGQzoKghjyb8boMy31uebcjLc67AR4VbRCMEZMTLQAy0srhDv394mw//h3+8EVWYC
w3zhs8DA9cFv7wJlNL6Tasvf0iL6Q4GO3RkFQP3TevWrxiTYOEeUOCNaS++eIA1VPQ02DpTPCXPC
Wnx5/3S4es4Eg5Du9WEf+foyC999+jc6l52+b/9bIcer+3iYwBfYbLTxC5hY4QM60lZaWw4+Dl+9
jZKrTxMfVLlLu++WfMTmjiN53ymoQRw8ip4l0PTZ2lMc16KLoBlvndPUd7xP25vr6pkgS5Sdb/Ca
Kfpglg9HX0C8LQWYWdmjD+Bmb80JgxjgyooCDez4aM5fYlkovXQoV8JJS9H/FuRmZDlUR5wbKhCM
n72KxNhPcd070s9GdXyuUuCgeQL6Og9QxewBmD7RF29vhsqOxjf2D4sSHw5NlNHEFC7r6VnGqnCZ
kxaMq1g35clruximXysmIK9SigPNPpKntrvcJeivIPCBq2M3c9lzPBdQ54xZTzhA5PCXPDGj/tEJ
gsMLrsgKguO2HDRfy16NjL6kzN3uwjKIfgRgW23YesV005dan5w/Txc67SiVJpv8OB6flMiVQTlz
6ApWmcwHwHL9snsN0C16a5F9UgPUcd23aThAihUWsi7wvyx5Z8cgO/LOt1MCDPCtH3zH3tRXTSL/
rIoYRH2rL2EJQLZqRJUxqTXutzkmECYYUa6dUsEIXaeZwLPPt3u1qHaNOE5eN3Ss/qIwZ2vsG6yl
X6Plehnf3xxeyu8Oh3QRQQhQwJDpA6+Oqtq53WR3O2s7oXWeWSrYWddE7QCkbOH+9hcqq5FblSaq
sM/GJAaOIAwOo94RrdC6/FmFs2/NepETCEXPZALG8j3oBdSsJP1WkMVk9CTl4I3wJ/xm6dtT9O2c
vWu2+pjXhQlayT6CNycSDS14RIPfTN8tPu5WfUSlBVIBhgyngxYzsPSRSUXVSisVsGYUfY//BDnv
MKMUfXXZnvC1pagfnzer6S9z3VNchThoZVHwj3ugmWf/0vHRNPjRRIw0uSM7TdNbAUzlcMmUNnZ4
b1oORSvDhfgmPNhYPAzEmhCGGLQo0II7esD0oT4qrCx/pyQs1zI3ExGdRVxDcQnn8aGzW0WUBF/I
tfKh41WV3msIbLAqNFCcCOuv/eLlwmPmaDthcRseDFsZRaI0xx4gXD5rZ5ZcFiXLkZpQzsVXi4Zs
zok9GEuyJE72ypcavJwRn5JVRgtLgyZuttrUFipXFtMn39ghpqKQsTyjry4dzdWyMvo0bH5fRZa2
sfcx5/QvXZOXIUkLYnF1TrEP0dk7D4lF/817Ps8c6PyEE3m/Bg4aUmRJSRxM0Hib19na7PmvitBC
RPEXi5JTzuqHkAxzEX3RuEp1mLqrHTqnM/kqqW5NQzGSLE3hxqME2mX0qk9jHrMuQypx3/g9doxU
ou6DxsT5xm+mo5w8o7urSdxFHXOB1Zbeh0NydmbiE0BaBaF2ilgSPA3gvTpPhi/RppUY7HiOtbEA
vT0V8GhGZZoWIOBnm2TiJEvhMYft3xY8bBhAx7D2jGQSdq2OFBXNMIZDB71rRy+leqs+pxqfcxDl
bKWtwBu6shzseFSZPRiNl+4js+k/7VhvWIZ2YbyRhKBRdOD2HGqsRtsqtts8YIgqYyv72cokjY8I
Dokh+BDsQ4GF70aBF3ufpBv4huWCI+hzI4tUjBQEAfrqJO15g+CwPLvAX3pRihFDQy6Ly/bXExyj
kZ5SdPhoaSM0+xEzHQzT1qU2y+rN99BmezgC66R+7bgwFjyxnpK8rkMju11CizEOqfUpYO0xf0Si
zIp0d5kyQKQS3wmrhTzt7gRZGTiJ0MKUwm2XBJx/Ia0bt3tErVHhYxkNEektanXyFt9wUAaauzCR
l7DXd5Gl1qiF1RBXusg9RHMj9xBG1uwEHDQ9u0e5FPjpAhFFTA1CO2Bi9BhL5lZ7Kaho62chwVQo
kRHOxeuft829bN9uuLRKq+H78TZl7vVCTp3i/UKmM0XUC8vPUiDUbkshRwlRqVP+cY4kslld7byY
4x+ehDcGVHvxJ+6nNH6umf5K5pgMTL5hhJnDm6A88aBtvqCHzFoNEune6zhz0w5COtsQYiPgYn8O
A8Y4/07I24pygRuRYI3BWEmgBwS826XNcelefkI/gcPEsEjohDuhO9c9IGPmpaInS1OUH1Nf04m/
gH85YtAynyJSHZB4iHN+Fam2pU9QaPDHvKMLyDY+Ylc50ZQrZ9IOLw+w/QzM9JG0nXJe5jD9tNZa
TxaZ7OF1ThzxN2r2/26SzQP1SsrQglXYgwRkXfUe204M2fy3VXXOvnT9KsWBKBc2i6yfDstdPYHW
fVN3gzVLBICvOBv0j/eRg2jYWs9DduyKm42MPnlDmbne7v32oXeFdzBj5gNZtODr4rR6PoNGt/13
Zed6N4xw0DVXDrqEJoc663Ga+Slc+/DCmsZThUe/rcNhlnr+fgRBO4W65IYDcPHGCbWWvEzWFXz8
nD3lqOCUCkC1EHcCbb60KD1Vap8kIK5qaS5p+IVP6LbkWJtd8HV6wGGdD2KE8zi6Hu16vjh1RpRi
Q7mPXJ7qf+7tXsYfZg2WzcBdcaOxV4FPvBAXU4GvNnclGKIvAFmVo67Wou61ldEvSvASIK7uShqa
5uh1JGSd/2mZQWH0nwEfF6dN+4FcIkpeInN3kOEIuANTRoo2E3C7RUP6WkhX7cTc8VWJFmOXjEuD
I40HefWcEccHoYvtaWAaJq81x6R9xR38HBuHWI+xuxiahq3koWjiAG1eS3Wo2S9bFywB767Mf5kz
QT1Yd7Ww5qsYychqOf5jEKviCJUz0wvJ6FtDQ9HJ8RLYWjeaLXCaqZHO78z1yyg2Jso0q/vcsO4G
XVDnkpcs1qByTJCReeQjoOIn45v8UfZ7JZPVEJkc/trArCme6VAor2WB5Gh8AvL/KVYTQK1AbaT+
DSPiyZYRJjhS9Ip2M5aYw5sEwbM7setu3qdV4vCPO7PgnPy4XWzIUR5Pqgwz+zoehnnJTf+ceErF
XkAKmUthls6TMNi1r/tXd0JJNyM87sX4093EFAP8hzcQIXYDhKxCNYqN5QAh+21mQdAliJqUdift
mWE5lf5EvCOg3Y7SwV9Wk2EmeSyYub5wVoc+eB9DtgQLoR5uxWTXIjwzlYD00um2z3sRkSXBfgJF
7Zg7iBNXa3zzI/kInM2fkYi9oyzx6ZQx8Rzu5U0CmUVJdeU9ZYmvI5mHubVajBHcav3Sd6AYncQR
UzmzSfxP8FjhQA0mRemCFtT6sWiWPuaymA+th1UTWurvrCED0JR2eaY8reKsH5KGm0KXCGNk5llO
T5vahBdCwEot/cB4a4wHJwC6jjHOVf0RcPD2o3mkZw6RtPWMlFnsEOHy1WnJPD3HJH+MBvZzUrom
rpxC+HV450cTJR30ddqrP56VXCqrqBSecQhK/ioBrO942kPz2KWL6VZ6oBjOxwedscWzRga+++FH
V/31+r0Gciuayb4S6lNgRAcQ/tWD3KNYXj8/pUUnfQl3LJTeK8hJG9LxUJ2vA8qauV+jGxsa+2Uq
55nwCTZHwVZX1cS60WBRJ/WijjJy2clXZsRcKlDuN2UwK+7swSvAQxUmX4v6SJGGBeWPtFFCnJDI
XWY3sTDOoBJ1KM+L1f2tgowYVmsvupryoDZ9DyxMGryPTlaeZWajFrNUkToLGlGhC6AwB2xFYRjE
LMmw3c+PeVZCR59h6GY1fgvCmitW9MhfZX87TWEkgRp1EyhObNehZ+vHwGcHzoVpBn+1jmOolj7t
3JZKY3rRyt4UIg68mixnVnbSmKEi7T8DfZVEdOJuRw7bbamkbrql9VNzoUu1gwg9qzE0H6fj1gdh
Y8B8yI7IdSdB34Yw354OX/iaCU8BYTB8lWbY8z0ijZU9YqrQw+c1N8V9eyHux9MqaqUYSU5144XM
5MUjWwzDqfapfFhEbmGe8e5AI7XhC5DEO4rYTolDwbUHjMnrNcS2nQOWfosYsSbx2bFoFzXoENUq
K4xa3fhycWzIN3pnZwS0uM2FwSlwlM2vWlggmmQdHJR4NgZudU/d1Wlnir+NqkAfbdvVXMTWuZD/
14YhFbVWGULAbxB5H4AiI700OtPpVMjJXA6EoO1uskFpP9i6oYXMRDVgaClQHtL6ksA/XWlYaUsR
sV0fXckjt3so1DSG6UKQiZcmV/YqXKZuEWxHHBXlUr6TFoL7qGdO7+dNHYufKgMonvOodCRUtwyR
n7oy25RtgWxSWtTrLfr0AaFA8+RL1bxehsyRvW+xhfsuaXXXy+FRyU3av4JyQFbRFfnQ77HRDels
ypPyvGT/osN9B5kB0iT6de5+kOF2yETUFZUVaZi3VUVZNOhtMVJPoSchLyEBnm8voL71U3PDur8i
TqzepdglcG2ZK6+ssXUgJPJZU9ttU/Y6nM0jsKbjQffrO/iAtVD/wSpo/PoaGD9ZH/ioEyPeVqw9
ueJOjS+5ILWqzLDuWWtfRV0j9w6DSDW60NOYbYOCMP3F3nWFzvopXlszHGgp8yAYuu82ymyC/7xY
fASShlaiKKXrZzF6eso5MScpoe4vvEmqBeyHj1A1nbDyGMm93/VL20PYGRyYORmtn5yoKWUYg8xP
K5Y1ERTeAvM4DFoZVmah6NlP6UaSny50om0/oV/GqrFE5E/Khiw7ZpUdCXuHLc1wc1YJunrteJMp
DNfgQHcPD5yo3XVNXFYNVpzd5hDzZqVqH/52tLctCBefqr4aAEId214nXxRPy6NH11RJ75Pp4taa
mzyxRjUvqhnRg5jHPEdnd8CgaADpWqwJ3/h7KKT0lXBZdDf+C+gLhmEUx9VYk3G/iCRWfXmQWrF3
Hit31gVzmQMeshZL7drPMacCiAKOOhFM4c+pM4k5qQbb6nHFdIfUANXpFSBApY7tpUx3o4pzvL1F
EFDpPaQECWtQfsjanq2MZbpS3McipqMmC6wrL7wQhl68V/0OOqsywiNR+lyf/47Q1+U3v6r4UXJh
mXIe07Ls0bXPISQkJl8D5z+8zulmT3woMizJAdqgfHjSF1rhka6HOwpNGxN10+fT2G4wI45f5KNz
K+4XxJnwzv2mfOUBEaQg+BY4Jo/KYlEM4X8/gI9Ai6VlQF1rP0zeLq14QuJS30xULpGIuVsohspM
h4IJTqE2nkRoll4F/Bv0u/goSwl9EU1rCyoSU3XrCqE+ElCAG4/A6+Smh2n8I88Pmx265vzKEXHZ
5H5SdbiaYp7hyAfjwg8Kj2Fuaup00Q4acK3/1QzAVXqVAr/DPlbsI4WOaHCCYGr0Lp6f5wfOc2I7
sdI76Fzah+NsA8cKerDpDD3GN3ucjBo5L6FDhIGjnR4rzQOqmk0AyZ1+GzFE+bZWmBQ3GNYXFGU3
BYgvvdjAhYMQuGF0hl0bjPZKZUf+juvitZw7SeLSHCmYm2uHoexSBreJSeCjH9iO8jrDMkPi5NXO
XtZT3167tqiH6wck+6lhzMyQusJVZ7v3wp+EtLJZ0McGth66Aakx55PO10aPxxXHUa9QwWBxDO89
d8D0ji5r/qsLOMKaT0O+Y5ZUJpKK+mU6wNhlAovpXPrF43oZoaDdBK8FJkdT1RXK5P/258cgOp1N
t1IISO1zXkMzboBgUcVq2u/vSDTliDJbuES5QCoA1fpoZT5qjAuf2H6GN4T45TJf1/5p/n0ujRcM
d5VuxKFPe0/A7vApWMWlSqTgtISiMKbRxFnnSVlIspqyZQNd0e5m6VKVgUXKgsGxCCWKVdb56Qgu
KQOpl+ogCoLRktWm02VqhLDUlcXald6LwdYXGxXS5jozbLIG2GUqpe36mbYYo7ecv7dUchWmJjlg
JSMVi6aSz5BuKdm5caX6SVyfUmT8wYNuv1WWylg5rm9necjxbhS2a+m3ZzUPnw8ij6BMy5AQ/hOd
RrgRXUVld5yyU9tjAOu6kxx2II55gaRXbGkt1z1S5NpZGF5+sODF0ubzCaKRGwEpTUABjsE2W0v9
cHQ78QWA98cKxRftUZVLryXDDGv9lypybHwSRirvgT75qfSTG3he7c3Nbk2iozLbH+R9gQrCFDZV
7CWLRWlv7okKDL9ITBnp7tPDtfOkLXDtTzmvD561HqdqwD0MrhKqSGI759bZVz4/sK2O8cTO9JSc
C4U+AqV4a5EU+13halH5aYXBjk3PXbTqC4x3qfE0irM3tE8H4HJqeZyM2AuEzeHnB+5sZv+boAc/
CmaFh2Xkd68QX5U4KHQLNUou3AgbQx3nnnwkfX7yxgw64ZULsVbIpJP7wAoIbpKS23eip5vHbVE3
7pAaefuVHxUbclQ74A6AooDk6QINwPtfPhLD+3yAeR8f6mXczCNSv9lOxNZC6+2f90YnKGO6RBOd
QPKCqKT9HWlQXT0aEsx2U+iFHjL+BE+uKk8ot5AJFEAx0yE81/WrXVlRPDZIj78jozitZQK118GQ
NY5xQPebrDtGl8SG3xFcfp1Z3YbnwdQVyT+K0bQOZuevBZj/AZ07WAkQp23O03MefRaAaK6rv8pw
34K0ZMNx1KcwpDSHWwG6Ol3l3ZWLl+vJNg65B+6GiRD14HPbORfxNXsA8jhgjL2FUeA6CZZk7Ek4
yTM1hQFNDXv20xTBFlYdzDjZQtQkwK+Bvd18R1moZ5G9VCGcgUiGefVrFp068I0zBtYBSAxP1Yg4
0nkn+P+0DAMyYGSQrwJsOlWPHb8R/leGRiMEI7DI2CBk18/YFRh3xteiSZpwrVYhkipGLXuearFi
LukOzNzHqO/C2zQjp+1RjpIktBX+X7qNgkkY783rLbvAqPlJyuTLb35hiLD7Z9ANSgd61TBd6xo3
Nx3zcsyu+2eHiTj5TBYiZST1GGxDfZzvpCDEFQ+2aGmeqNGmesxyHfDr/kYyC5omMujVOUbEwCLI
FlXuzLAnzi3yLardf+SjIECtoOZwEPqvyDrtzwkNK0R+i+aXnAF7aXrqB7D9CMPXbDoXERNAKYWO
BuQByASyTgoBvUjS28lzY8YQC2kiXFw20YmBidRhB6QioBgDCK0UQlTXIzaBuiOc8fNvnbgq+TJR
WYM4xTKmXZYiWyCU9sHR1xw3wDvdq0cjUI3Ed4avj2U7ElELyObNSzpoGltpRakiXGQefWfPS3ve
3XeYRVqDlrTSN/6SY2nXXU54k85WWx/odtvpwb+RKfs1ROls0YQypZmXuO01COyZ8qo5XxGyuRa7
TBNr2KTZJ+yxBkLMY7pTD19ABAwBLWqLz0xbvIpXkz9uSPh12K251SvjZ/i4jx5VxD1mmUNDyXPH
U465EbGZqq6bsmZeMYX7uWmBLMaj4LSqvegKPYyufkeLPPRW3wo8mgqkG+PEa/Nldcg753P/i9mE
Zr+EvjfMQKuqT8r4h3kNBvPq7aqQSBoB9r2+YiHjTwhYvMDSnmvAEnt0f6XAg7aeqNhwH8Es+dds
WSi6nLDVFgre2EpED9fCnVFyZ7FoQ7ovIXJfOisCifRA3GbCTTzE/zu/68ICzJA2dqsPm5kn6TSY
gD4sCRZpy50t303pGCOTzJuSSrCBpHTXUc8ZAWCwFfYwntYR2GihU8H6HoF3upv2nBA6B7Ncyxwt
nPeYeZ/oVnfMelx2o1km9npEtlHrl/G2nQy7jM95iZr7KX1wBf2MxzthVfWFjJ5RwNES1juuhpzg
Aq3FgY7DUxze9fwk4Hvsu63Que8TqC4d2aLJWTXgjy728Cbc/aGYk60rZeETx8TrBZE8MLuZutY1
QGBdz6bfqZJ3kqzxi7jpS44X4ovj0pu+G5ZeTlaMJOd9GCv47wY28oVpxi97NzYQ7dlFSMpYMt/d
U6DNdncsW1duBecNaL4mAGQLaWS4RMUj0BFsKDNxh6Lp5iCeigR8rqNgTZqyjBekKLPppp+nnOmT
2TEEnNbpM+Q5gC+hAY9KxSgGb3S8sg+xTUYNUzTqUiKAlxH0Rrzb27wsKhR+3gYTTeSwj5/uvGi/
BRGvEoLdENnjQN5CwgOnRpauDSapYgQLIF27Gd5l1HNEvkJgP2Fbc5AmldPRaIEkWKvsJEeNuJnP
yulKpQFNdMNJz+2iGRlb6Hz/nlOJ7PIdvNeUJDwuEqxaWD3LeXUQT2ZQsebkHGdq7FMhbqRcwzqN
hbSeErP5PyhwpVjg4OaU9BMwftlAc73Q9UQ8CTOrq9XkDO4h0oadqsltd2xM5qA7NBRM9xTEeUV6
4q5MRjgdN0Wb9eutgXgV/PXKNAJPqytfXBm9dw5R58AYTOsNcb1KWqad9ZQWbiDHZbNwndE30rb1
Lv/lLBlCxTnjKBnegebDG78byfzkYEwhySlpBHG7xbRSoKLsbnI3VMuMQMAHjV7Pas5X1WfyCeW2
mIgN3k2UbQaitI2DaOw9GkBfr49ak5Cj12JZJ4RA5mXvUFPKHvy1aM2zX4zJvKArm88avdf/u7g4
ocyuQU9zWEzAlfPsCzDkCZDQ8VuBhmUtXdrKkFWWmR/GqOXK9cIb+FSzl9y6J/hmNDnkIW8uOD8m
4EnqBsHgguRo/N5OKwVOofBiC7RoshLD9NWVqx7npc5sGFK+uKMPc+Gvypt913gJwdDT2Yiy/Ygj
faCv4p+UOng4dS/IYYOcpDakrn9yyUv83TUAMCUTZaYBzcJKqmt25Zfv3jqN/UaH9La2Xo2RCrSs
r5wkfg8FR+p7OISDKoYJssd4QwbTpyg06cZNdNs5gU+i/DiVmA303t1Tux5AjRJbbbjByoJ5WyG4
e1JnbHRwLuSgIkaTQqybVgTv1OkE2cb8IbuO6DV54PG5Oj9HlgrkemJv4rKtdwc7Hh/rKHxvpjI6
7abhClUQQB/EY9Xy6qs0VuxYnTEgMBfAPtLGhZJNREDurxLHODfgIpPphieuVhhl6EDA6oZcO1Zq
6ZtSyxXZ+HxPQJCJysXybo/1C2CEBkEus+1eg3r20Qe7XUxE4e5Fl+uKZwoUioIGPMYa3nyqnYoo
6rI+E8aWur7sa6hGkI+D8T3TCdTAnMl+e24L7yyirzH9b2FIDqMjLHw+uKCcB92T12oHGVaFejC6
ug+TmdTaQdQC7RI5G08x8zkJXYFRPL0TWk8+Wa+ucmSfcsl3Y1m3aExxwL2Ew52jUlVSLVJajtZw
nZeSCmkhTJiiY4X5AoZ3+dtRdhtnCoOZ/3azH1ewHygb3UFmpRP4nvfXWowodQNCBOkAtJL1zE6U
rUu751BMVOD0Qkv0VDgaKdMIbfPiVjZoukJiTTAyJYjmpnrvu289I1cnZJKOy4PRG+CqpKW0Mit7
sNKCShEUCOqNZ/vcVBMsOunVqYb39qPM+yP4VyUudjDNH0kRPTVQxwfqOw+VFxAE+8X5NlJ82jF/
s7TbFkzOZk6Pwe/cVdHRvo4mu3OyP2yT4YcEQCYolpZiMWI8/3m84Ad6Nev7iOb5oA4NHmDEBSVn
X9aQC7qFiGR2EB5idzf64KUcQeyepezhTIKL45H9feZLNhuiM6rR+M3QDD7qT5WtUSmsP4lNsIsL
awsfFWSTXGZa8jCQFWT05msabsLTLdJIvhJ2DwKr2BWkfKP8BBZV6rfpGgfW75DHdsFehTX7hTi8
MbJF3YINtb4mM9tN69sy8+q+VRKQsmLi8kOTFarZagguM2HT3YJcjLez/nLIGww6SxLKZpWgq0Wv
iccgIu+bZS/35pMHlCBNi8HtEDWYctF1EE2Ojdx1lc4Q2emgYyd07lljRq3QSSr20kVGCsqnNDKT
9uJcvLezLq5HSpGTtl/1MfaVujI5iUz8+jKxuLhnC6LpQrj+YfSiTPfB8DZfxebj2v1HY+5LAe/c
AMxnIM1ULQ3WUNXdXPMSWImSGcDgBB9x4bmmEEizzBzYz2pMFqrkVZAVPo3maj7JxZjZCWBKMh4A
0+cry+V7vTQGj8ObH+kNq1X+6nEmy3ZBL89EYHxOzp9H0Haa2Xp3+pS4QOEtc4mewbFckqe4PGvu
koLpA1v+heyk1EWQGLKe9eMiIICcq8UVtaUAd4DrE06KROD4PS+TdWhmXTAg1YBEMUnwrG//YzCb
tnehP6UZw3c0ssAJquMa7KKAwkSXKWnT7hX4ubzyFfSiSZRDgFLGQ8oqL8j+bWRQ2tLVgIiQM3pz
Svmft/Bfww0WcwFFmAeAN0i+OKmLzhAjYFum9RL95gK6oVI3UeG4oAlrVjaVx44Z8lMFpA/uAHjX
OeN1Q6RntEmvfidzKA2J1Xs8b6WrK+U0WJOgIFaYBjZGbV23dATV5w3IRxrf6/MUkktG66VDoL6u
2b/3SXHqoxDK7+XRYiY6c0r0PRgeI9iF4/7NCbx4PNPfoWMkAXZwZy9J7XhE3/1x7B06rozfP9Hg
n9ZEMXYQ4B//Fuc9h7ZLFAfd7gC8w3nqh2sCegxdpA7QwsPyc0UIosaUyGe44I4jX7lMwuG1LyZT
Vc9bWyQTHZOoCrjr9NN0U6lfxMYqtkrlOtxHgqhdx7uA8LL1sH/FZWRBXAJceXybzhjlk/VDkdY0
oS/7OlGXG3Yn4UK4/Th9dQ4KaxJSnUYdG33Lc1cR4NBzncrtm7RafOzIL/ucw1GPYzSgCSTF7bqX
462ndqpCwoH/1wH0CJ6tnc6qF+K7fPAEPbP/vMtshEsnYp0KhoXlBsVnkI4016/VezAfjdNnHMun
DUKf0WIQBucb9dV9vh8wTzsngO43Em85389vzRh0G6IlrxJJMVXkutK4xKNOFObi7ekxRM0ROr6X
VjHeuXLILoWT7dyruCipHiwWEhEuYDNmnQqU+lNprG7VKmA5o5C3xax4g943San6yBc/vyB+ufvZ
GyE6XK2jokDAifkCnlmlY8cpYvQv74py/pDMN7tieUHhyDDMRHlCCRqo6qx+8vzFTLMJrlsGMeY6
CMkMQgu5Mjm/2kGrrf00BfgeB/BVDtDP3Wf1Kx0NaHmd2M1sroyVz8R+gyUB/IwbEcBBDhIxjoZ+
fRY/aAZxsrttvL1rPbBTCBG8SYY84q3q+BTrVZ64J1OaoPyDU/f7/l4DVDUub8LXEW0N9OHKv2tG
Kq7gCbqY+qQB2zA319LXIImywdZpu1O6yNvyIVHg7P49WPWXEiypuEXT4mSM6xVnK7Sy064iSSYQ
bXoag5F/j3u1JdJtziWNDOE3OFZXeQVQ97ClDLBqU+LS8cOWUIkzw8AG5LSbrOQ5C8JnuveH6lRk
ewcw1kFgAzgEOpyu6H6hLyp3Ih7srRPzGKXf7AGCUhm+B9sGC2ZpsaXml9tWPMiBTAkJzutiDRrW
AxSVqnA0mkUcMtNg6MCV9+TTautd8f26lJ7cYUgbpd7hqqiSKUIOqvO2UlnQlJM93BfG32ziNX0C
/0JEZd95SRBP6a6rBFK0pzcZjGZshPhpMnidKha2/7NYG28CU1zh1yViQsK/Tr/wrnA3Q3KQhm+J
26xFUbQeQjeRSu5JKo33KHHimeb+A9icnrkpl0NMG51m0khPOwcIIVvYvK0dpVZnlJUi1+MZORP5
oTT2TkieFwTla8hvpGSiHp4TH1EJ98VtgRnxHJWYdz3t+kbBFYDMvGX/aRCbkNNH9Gqv1jc2465J
Lswj5tMPlL+Ovo+qcLakK0uCBizzRiMmwFXQjknIxWu3q9vduIn5/x8OP6ACPGHyZU48f5G8htzv
Pmf7Osc4eL/JCdD04wNXg8WWfseYUlEHqIBW2dU3kZHsej/SR71Si+ZZ7istSSBXYaG1PKRDaFXw
/SpOYnOr8oXl16CMgbzQGzKCYC34OJ2FJU3wLKZu4uy8aJH1itnnUxtr5SBTZ6yH6j0nrDUCzDuQ
kRNW3ZIkjMUIDQS4jd8N1jCUyt9uVogixGel+JArs7zFnnuwYmDC8PccN/I6MFsJ7QtY8oxF/gH4
rBhABATxlTo7ayHoLs8AJGr1oaHsPSH8RWzK2RGblmNK+WJp8ysd51cdpAJEkGvNf7mVs1lVvxgb
ipzRvKYssEsuz+EqkpvvBqYRGSWJqtV+gvsTIEZSLgMAUHWwE/wUuctsdSpabjAW59zPqD0yZG5N
X+WuLHYM6ReP4k+G+FegZC5YGnyLZSWpqdPL98ufslPF+pqLTEzf6vDWmi8X4n6I8BFCsDSRztZ6
jIgxF+3c1TgcdkIAIDes/aX848TwZlw62YLda5aOVwktTp1i3hJh8rjldxtNbC6qo792BCx479Jg
qLMM9jRIa/uOgEOrbf19qUqTT3gcZ17sM0SLD0NkFiFsvDDsGGFFu2u9hABGC5P7h3pqN3kOOJuu
X2hp0QDRgnaW1RUu2hYjTi+d3jk0UmFxG6eYZyC/RC5p5Oi0fDARA9aqiShYuuZ6yv+HQtzgnC0l
AHzCkvJGRq2JWPRpk4nH/+uJ8D7xf0rjAWZnGgAbq4nzvp6d2FXeEizKz/fwiKAsCr+YJdgBPNyt
pR/8tanDYHqGi1J4BbfscKAqnxeaQzpL2QE276N2aaXrk3rHQVM3s6cuJ5s/H5zuIT3dZCEHn484
lU99U9rlS0mJVp5mzq6ah7+2EBGisLIT5D1c/WO8Qa+zj3YTXP3hEvNb3QLFj+lyqunQkBgBDnAn
5MmZqyuqTUGKgHtsm1ovGu0yfzJNq9J8nVHrBM8GbMPmcQ6NymSzuWqrii5RC765ZPyeO+z2u8rG
M4f/6CncL+f8WaiLzstQKK/nxAZmd4TQNHUaN0tN6cPSoDbJ8sZ0eZTPCQF8D/ZPXR9qaynvtfq4
ivqJ6WZa/HVlOtmFP295y5cxRLFhp2rGUaKCIA4TRoVAByaJR4ngsrQ3m5ohTC1I/9RVf1OJus1a
3rW73/VxAPfHDj5AqtbSGbB+o5kUB93nWbw1rWILeKjpBdbZvxjKOa6E+FPz+Ipu7XK2vbiGb+tO
KyWIl3LHZTd4ayTsQA97OIqMs1c2TQdTF6USWBKhbNN6AxaYyyDefwuQKzO11sG+Ae4ul9zBDNU5
WNc4FW5o5ORBNx9qUKickuV0k+an5VvzFCwb4DQZScVVWLFjtD51G1npF27QlRNlZxbST7K93zOS
zThJK/JVXEh0Fxl9giFTD2sK65X3tvO66NfPc8YkICgOQ9ixT0VGobuYouaxCvt1ggZMYgpe5PBm
viIfwdAHNQHNYrfRTa0En93gW1zMD5F8rU7s//b2W9Csao4Wag090uu3fc2hVWu3C7pV9jLtySXw
hErTn+hti3BbIH96YkNFhqlD6Psn6XJoNqJfr0aiHRet/dehclfHVt4S7mbgQkMM9w8SbiZjybpC
OG3gSYTMGYPi5TXnU7JNDm0LMAvEXbQ6HJmUUnZVpgR0f52j4fqjKwNJP9eRWmDe0B0I/R3fT+dY
7d0a753fDsuMt/OkkfzRpsi4NptQA7/uemuSRLCqSmLHEZ8B+FYFeVyTgDoAz56RwttueAjIEbGc
VSVxt6csPoZXvvpA/jnfsrrCZzTUfRwYCknSenXqxsTJesKtpYi72HmTjoNfTldXA5XTpO+N7Hk7
2CQaYtDn1wokS7Vj+nTvEMRDa3pv/mYUt/tha8jEizetSCGR4EmLlW4Vy6b7nuAV9R/GDWlnJyoi
56PDziXnrT89qpvX+RAGS1q4Ud3fTk2bofbVTMdfkqMX7WTRzaWlw564/3FFZPCZJiVEJu5xWh04
qyZRkKwUsqkk3k/uoa9bNJdRAys1jn5O2TrEPvwflt7Q4Cu5HN8wNvxj+k/LVYUH9bfeP3m2OKat
zqZymPruRgK5eW1/wkkjUb5aGquTbAZHp7y1xR45XX7lxnQRosDd2TDjWAli2oWdPImVVONoe8II
oBIYaXMoQCYlq0mzGDjq6xVtP/5Jequ5USC0UR+kS+5zm9PzZTmYvvyXguJ3BNO6IGHVnCL2w3sR
nfZr9Db7ZW4JN1AiQA4kQZTc49EGYp2Xdc2crvWNp/3T6X5vELLMGZ2Qjv/MvqTuFslSUiuxc3mG
87oc13zgVCWOwMNsKnZhIMdeQJx0hbAMi67Gzmqx9EwP5JenMbAe6suEq83pHcvl3XKkwTb/fGFm
BE2HjYY/8NMnZGQ8MswxTrsXWtLZg4i0Yukmj2rynGBuykA7NmdneQfgkLIQ2jL6evVtw3oFM2AR
4CwJZo2uxoelrcwy4t66/c9RIRDQJZoQbf33OopLYavskEsaoo48u79jmvQ4wS3Ks6/tLQPZgTjM
ZwTlRbXMX5msnKMnKf1uqcTDPgUFKwlYXPxuEqXqjuDkh5PIrUw/Xf/GyyfGySp1mtfpjEp5dcZ0
XdTTf92TWn8HvP6rDzRTvoY/wbaas9j3q7G2UkEFn1Eo5SQ49HAFemEI03PYJpoHfOu1nAcaVNBh
/fDVJxuKOsb3fvC9JC7esemF7oaX448qu/VaYxclO7t0TkESwYfGwhMY4U/CeVNnw26Rg/HryqQ1
NWpKfoP/j0yCVQaOEG+dlK6wOJzphgR40/ggeFV4YWDvmWLl3tmO8wB+MBhquEHyfuC7Sv5GfyWp
SWaq8CEUk7jU1XRtOG9aJUeudCUb+Cs5ICBWdUV+69O2YlWVcExyFXdsO3ZdIZj7m7Te4YPF2PHL
3DcXf/88E6Lvwr7CTfmuZlrNItb//jpXeXyQsIiPOULh7jqZ66XyCta1CBpV7BRaSPJ38WZko7Dh
GLGF28Tr0bqq6pAPjXkz5oHzTid2KihDqT+LM/Ue/yjOoHhDcCumxbLVjsSE4a6j9f4TCTfbpLw/
P9zlcGNEt+OJQjzsFRLV5h+ozBbMw9esxev5qCEqe/PZ42dvXvQNdEBk2nr3s9jSSS+6owC2rmoH
vePpZa6+jXO58accoCKa0Q4Pp/C22+uUMqbBxj9wnKgrH5sG7Uwx9QQYcQCNf8403q4eN9KkH2Bj
t+HPOqpgv4lFDBBFuwru00p3mGqB1956QdQ1dehCRvqAIXGTgSBUoHImbQokSzYyghlySUosrlXL
RjVzWZ02mieP1p6Wm54ulhjq04YKHSGMsP2HYtmVzj4rxpZ+1GGfJklR3wayyG68Akcg2O5mrwdP
TzgBknYCXTqg8N3J81l9lW+n9+BqCiw2xpmyPkxgCC/8R5qVHJyudUzIjOUwk9h6wb1OI4XybjFj
LxNh3fJR6ylgPY6tBPKmR2afxa03hkvHrNJHmw4REbyyi/2NG9kFoXnbQRT1VfGjnfSxNMHq0ruQ
MWfhnf8CewyzdzLSf1OVtw86PB2Vr7BbWoFAqlaV9hyUowD3zHy4JeYmstP1CCK6auLMUi0ALOCF
jUg0MKaoeh7Ot9nn0BIPqyRTluzgfFdrtG0kuggoicfnUttNxUCLs28NJ5adBhlaLvoZyUrG+RiK
BbJl9IbBoCXYhwY3HJY5/ZEx17AbDlVGU3hijP6D3cxTZR1VC1fMGi56OwKzvb7j5sP/Nb8dpVTy
ba5V7lqMeDOeAvP2WvyDrPj4hiChJdeBACeY99yi0nkhX0oM1BIIk7rzG/CF5SWj+kaDb+sc38bR
rNsgmP0UIT7Wrelerk/htAR2iSYxavIl0pDrkKbOue7nPNsoQIessG/uvBmbBq97TtJylxnTIGt5
PiJk7egJVsYrOFU/rnXdCPDEv5nmkvK9vpgNt7P45EwUBwC0b8/RrRDQeSBHuudJhQF5PKyT2L9I
NNH628xjWO2LoYnOGFKUnyV9fGhSRa7g84p2qGWdYU4wqMTrTufZdmAbEAJTUvJr9SWj9rUDDCm7
1qUlr+G7mwLfEvd+WFmFl24hbwTApfj4KH8NVGAHLCyTZ4uayM4cfNkWr+ACeO+dGaHCvtkMsWHA
GBQhDwYa9zGJzqHNOLX/9DRKK36goGqAjgq3t5MkcIUrhmy3fZPLFkByjCXxmbQPDzjzEvJ5054j
0ILicesTMKZ92+L3ucq3kHLZQbEiAkKkec3OREKT0p6NelHMat2RAVOzi6QLAgqpt0FfTsMNIo/2
wIgcSMLee1jTJjx/HzplSWN0jhMHE7SKVi0oBpt9mHZ0AyBKzzfLbIJwJbzTIUm1oVVZtGNomCDb
kSKcQCRAK78NCofJ/KRG1eyXSnKuZZC7BMa1e9qCqme54/KkNwnthDdWF6J5UVhlcqmmZKpWYfI2
WKp+a7C4TDCtUawvfnOZmBw9xY+FYKp94J+TIHQJWz2rJi+ZWWkWRqljGFPOTrV8lfb0+O/njlcQ
M3oMMR0Pyvaz3/sXqHIIFCPln6SKRVtGOObxY70Vol/ZyehFaPmENru1D8OoGcrLM1AgR1Va9GhD
IWVUJKFjf2JIUdIPep+372ZDvTbwdDUf1U/ASd+sNZDJXTdA19va+Klcfj1OglMhLfuAHTseu63h
gLnBUYd1MIj+13Kr5axX4f3vfsBQYX/+PRn0FaUntPyzHwM00J9BAKn7WGwZHeACRqENMbISw+uX
ZPo9HjoPANo7v0Ae9ejddRu6FQSbYLMUUtWgParRIyRJCvBhxoi+P294ML6LB7TmiRy4i1OeutBd
4Q14VbIVFM+byXBaQd4bVNSg9UfZQssANju/+tQ1IPCy/lOduxo9/HkGcuK2dLZOttffqMB15qt+
XHzreDso2MDV/HGXmdd2omQRPn94DIETTNiW5ceEtvULpgoD1iLExVPlK9/HIwN2HKyf+7inF3Sl
rLmyNR2ABBOj2o38K427rblYEN/QegwwemVTsLS+pJFHKUKDnaFm116MqSTeN9ApTqIXFETt244+
kGHYd6auzQsFitabbjPQcBciVwR+Bb0fPgAGAKI/2lRZ42xKkOM9WsXZprNAE4fkDPp/uNF/fn3m
PrTBI4I2LhuFTLMznOlbcablapcKUZVfFJ9UwAW3Nx8ZZnPg1P55tVXkp1mJ2LikIh1vzDhDPHsH
iTvArzgyKkYwP+1CF1HLw1dIT+5/RRzZwLYx/a9NCj/t4fPdR7I+fihrZbLT0op7wYJiMGeM7wbi
RCHSwODlDE//skKGYUlbLClxXzfofcpMhaizdE+cGkM5S+mYPmn7FZ6EHPq2N/gbaLBiYz/Ckixj
I0Db78kNs0lSnoIyHJDRiYu0FcfRqr3L1WUNEec6azOB8VSDLmtvDBF+kHsr8jE0bkrAPYgI6///
LkjQGr4ZWcQ500ICSnN2rWaEk7CESedTnrAUVSgBhT+IPUdjlhOIi1R5HBlZ3VCBYmc=
`protect end_protected
