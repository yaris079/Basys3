`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
RjTO7uGlW46CD+1ghMDk3IAwAeM6iB6Cv37shHugJyODHDcu4M/kFyeX1b3uW9QwFvmmLOMfufff
0+mFPegsDg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TCdJlMy81LiSQM13S+raTKskZjxRWNKKFSDalqoh2kIp2Bgf9yX1UO+/C4ZxJNPdUamQdXPIfY+x
E2O/+jl6u99TPPdOqrmyL8mYTlfeMBA2STjT84XEitJdLOuO0vkru3WGY3kmBUyBjCebcvHqpzAH
oRKxdmp2Bb+N7tUhhQs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lv6VYGUxXvT/a91M2WA/MQmnebG/3XhHt5mQMKMzGqOX+fKZj/ddSE8UCl6MSu1sDtVZgGG1GjKH
prYMYUvUXewexwueaNjkJgLn6gJZzGW9Z3D275q90BL9d54AYpbOdYYkVw7rkSM689mT+HTmwPyk
3pjNKXY8SjO7gNQjohyNfvGwdZp8w1gwEg5Vp01wW41XGM+WgTYr4hjIYsZ595OnlfjqiApGpPm5
25UAKf8GQJhHFvLOpKySbHi2J7mTAym7+P8nyMb93JWg1utbew3m1gBPEbps0KAz26R7sRvDtWvx
MrlATkUwXZg2Lc494ScfUvL66dKWSBgAsMyaeA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
v7AkG1QeOsPzwACZEWmzNtxMPK7DCKTzHpMr314HhlrdsvmeTQmys8Pd7bImEa09eLkQxnkAo+Qg
qLDph8GPUn3G8U337AFuhPjMepxrtWvjLfb5UXgGysXw/r4Y+Dfh6yqhKHqfUlWKvVbGv3PDPjvE
mMTPvc/0bs9XeDoht3w=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ENBotBUCYnCLpV65nlxe2Z3cGSyAkRSeQKoghbde7KSOXsG7mSMAb1KBMAYW5AhM7OQ8rj/DfRgN
+9+ePoIJCm4r+D4lUZz+aKyX2BNrc7W0SKgH+AAFxtKCWlLgaHeTIu61dI2lYJWbxHjBEdoVgojR
hwq9Z+alES3Lcfunlm9TRKdd3r62/lzmnrOmzn86cHYZWj5kemebRhauG9ThzT7xyhBmti57QIsf
gm6wz7bl418XQAH9qSL7/B6p8llVtWmGMomqNdsf+dAPZ3NdeP3xQ4pBxdeqU2I6T2DAltj0alg4
kcWGpDzP5riHONZ4IFmpqgcgUzB5qrkIC5YzBg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4848)
`protect data_block
UkJkhGwQF/XHARcU3F958O096ZUzihOSHOilLm7rZ9wE1shIGpYd/I2KKwIZzf6OeZTCbK6g2xzr
2JsbY2GnPwFg1WhDuET9B3hOVeH8VjpALjFIlDRUiB/GYA3R43ptUQqQiPLr92ozlmivdWtLsBNf
3TEk5iUTPQYxN9StnxPKfZNGdvxhIOOZUI50cIrl0YOMjAr4eiHk62R4FzmpjXB7W1SaY4U06/Xh
JDOIRCu4QtzuAmcOA6su8wttW6n6gTObkplltxJooH9U2Ap2aiTGaZW227Mjg8uSFlEjemR4jzNF
44GrhUSPhxme+lV3yZ61SNisdVwhmsgY2fNviGcisLqHGvDgkEBc4nyX60kGMZdt9sA74OzXu58F
0LSwwzeMHHiHMYdz5LtQHX1c9w+xMJv5RF5v0zCwz5tjQzQE+BPlifF+2bxZOFwW0KOO9KYYqRMA
LfuFXAn9bWtMImYGN8psgtbQ/3HX7VmFp/6fw+o2KmPPbhOfYwrrz0fORVINRC2d85CbRe104bzP
zuhy4gP2NNVIG9zQN+uyPjDKRYY8dBN4LboYeAk5sUEzAAx9dzNW/hDSGG4CNx+TNBkCrzDzq+kE
+WDrooB+PWQdsgyky8xp3gdH/3coB3EhjaDHUNGl5K9N/OMc+qSpPSjssZ1zQAnX9dXPTpBiY4rx
/B/qLQ7wUcb5qRBynDVgOursfPTZQou3qWYoe7X+dzGmPS9oHFhAuj7vKfJRxNBotsIxH4+fiEBM
ZLwMVnVxq6QWNjr68z1XNQbrLnrS5Gf49rYyuAVTqR0fqucy5bnzpNso/VrLJ+fcb/tbOgan2heQ
5CHbSvILwhzIx+OUozumgT7gLO25N8Rdvq7WNt0lGknUOF/lVVcKvrZF3x8my7g4jMGEf2p1bbu9
mYYRwjyRIPQ86nsi0O2Jo+eiAUe47C/kqvFrbY620sD1ZidmgfG6TfsXEeuli6ZJHLG2EuyLJSOs
z1pF+7lHi+adJ2CrfxiKn8dc1V/3+kKd3YV8ZYklOIQlBmV800z+i/UbcHqf2k4sO7rMVoNexn6Z
IofLDr7vIP3JiT0S3rMavNU6SiD3Se1hp8dU/lB3/YAc8Q7MvvQBLgzz92e0ZlD6qzt2Mnk1tCj+
SQBQz46AJq2u7+cNdEqjb1ASIDP75UNXr2dKNkEdxbMxcclNpitFhdGIAdyeWyHSrY0IqsZy94cS
YahTZEY8YZF67f+VZnARZTAmsXxNv2isnSwrxOz7pxAZxAIpLeOIGdR2CAdyPXJh8PSs4Sk9mTus
eLPbmY5kPlCu6ykery0Ha0hx5UhdKexmAbrL+OhTekOd1GKQCLpsZacjChFVQMtXYJbP9GQipHp+
KDjBI63Ded9VNF2OHKIKn2xatXdvNlxCAy4q3t42MZ27PcR3ldWkLJ99k3NY0ChAgx4fxsYwfUCc
8ZMEIOKaqeZeqyuBFQnaEIofvGXD2TbDeNKeSxLGmbcvHALwMSh2C44oeNDygAEB1CzmwX8BHFz1
mx1YGZWJDg0hEQZ0NANfoFK2HkUvN+nhkFTPrtYFn0TLXeEULEcGheM0bYnRFAkKzo3p1HuMvSoZ
Lgcq+fYGsxpIx0qXucqc5DoAmHMtN1fTevIhsbuNIY27qo1t0i3UA/ZbNNxPqtgqhONp+KSfC+hg
exvZk3zlybwZe2D0peunBp3+G20aNyXpw4I6f2PN1J1o7MD31PjS354D3QMVusmGqWYmhvv2/XZ7
kEvm/VZLFVXoJNpDSOSonKfB/iEwnxpZaxlX5VzGKQDUGnUJ7at7xb1KQpkV1kKovSUKxlQMw3Dc
yEsPQcKsVWEzPKNqC6jh9leA6n8E7nHlLR2R5W/j3ueBuzO0tx0jNjAlG0mVUWuPRK3SPmo+FKXh
RiETJPOsgshU0nEAt7iayNC1BHR9bWa0qeuhqodtiT1vJ6uReBmegfuMQ7luLMSxP9xukOAOBUXr
R+lAWiQ9+054hnQWb4jjNzpcrw11gBmAku+qJU8lniG6UXpTVUa8+Gf7sdKb4tgTqTsnPCiBnQWG
6oT+di/hWFLXSyzJMer98WjDzKCrr9j+MoBaOPv4FgytLL684yB0M9icLlGRYRpS1NzeQ1cfjR3o
7651jx/Yb/7iyRffdZLdalBViaBKX31CYBzOI8jM+GrA7FX7/AEcSq2nO8SS4TVdzmseKhhSNPdc
/Fd8mtcKoRC8szBwfSvcXdLp+zNSALKuE7GahDWxB0yweDGQCNGUahEGp1jbyINR65+ug6Mg6KfX
bP/vbrMX4JOp5sPUbZcMq0J//UxQ6hrbD4Ym0tnbdAQHyB9wLfSKqqS9Xa9M8CwLP0rSzWkvYQ7G
RRr6KKB+9DjtiOwMAhJ2atH/F0AYy6SupqMgFoUcCHD5r3IvdazG4iJS7jtfWt1n28dqcK6U4YKi
KZfeJ/96AG/tlzPX03/FcP3yPsVSCBtyEIRQ1gkRyeEX8ukbNeiYMRATvP+g3q2txDi7TmeE7WDS
aC8X0z7GxU+cppvYJo6L7NcJ3tnefPBfWyULpqMb23/ItTl9lhWBuwfpzFst5ddoa5tyU4uuS7YT
sV0uz7RmiE9Ta4nAl2ze0I6GnrTSu8SoBDretvAGEzx8tmT274XhUB79OLWgmH21NvPJp//Y7So3
QAPbiBJrRPiwoK+YB9fADy1fNo48Is1CuZu1Ow8G43tJ4wBqaymQzk5bL9tmVyoerxHwv1YlCHnC
buh0wApur+K9DnrWmUbb9lwwx4cEKpXqkFGpHBW0Iz966zM8dNEyp59UJlzRYGOuVk4+5K+9/XCP
L+wZrYx5MzTfdjjJySyGlB7xHqQc9EyWmBf+d9eajSO9wMCLaBa3G2SaiJog5BtjpAzkWdMjjOZt
06rtWIj/ahLSv1BQgutd+emSbn3Hncn/BqSUabqJUbDrOhvig1gWjRtGJRIE4LGAS5XL/htweHoe
cGQU5EKVF50dw5uKFMSPjXN3xRRWg/JnIHYbKVtWeUNkusbbMQuJaSL1kEPmklsdu86wgHmZgPxl
o1BnVYpvjThly+W/S6rdqMp9lOno0QyXW4EWNpJCBunmH4EoIU3j9lY/mefVaX8xQWsOlvu0mlQD
1ZxbUR0kVSTkbQnBo0zmbQSg87haa8i+1RFPBQjm2HceDxGfS8OlvBLj+EGayOGUeq/WUAvRSCto
0r2lPrk4btlcihUn3OnBrGEVI4cChaDvIED8/3vqLyZ5JEsFYnC1KLElegta8x1ZIm64Pfumnu9Y
Rx5f8BL2Y3fjGFgiw5MHKJXnN6SXaL6kkDD2WfyAHTyHAlixdlDUKk4QcvCvUm6DdgFAes3Eiysq
cylE095NhggDc1X19fTE4dalp8KgPf3knp9Bj+9kMTONP7Ze2QFUGw5kVzFwgIKnM5ZI7/Q/zkM9
YbpBOhUkcIXDPtgKbD1QrwikE9EnPW0RPkc/2YA0y8DYRDjtUj9VBuBzPD6Isq7iuTuQarmxcze7
B11Mwz8RFgOEUIUDGbL9veEkXMImi+zJpoIOW4kvp0SsB1XJ62PmrwsZ7dt2+ieleYQTHS8PQAXV
r5uT8BQKxFTQhRBdibNuS0ojz8eokZ6rBq9a/Lsgq8VoMBp4UWxvMHFclkzYPzuZl4bvOpuwe5Ej
IRrRt3sx7M6TdEHgbUso9UDzk2f6M9v5kvli5Fch88M7hoDv+fit9UybbWLz1syX4iI9qR8JJB0y
z1kGhfpCornp93biuCB6mSRrSGzpyrcjLVJmEcOo3+wDyPbYPxtIEJluYpJEzsNpxKMrQrwWlnUk
nG2zI7Jpd1iBoxZVV4EkSa8UA6raKVXBig1TpoJ9PzBUjPsRo0ExUL+DXl4+4WzJUDBxsg1TJAlY
yVpxKYaAj8r/YJyzfA6hdeTeszPl89zIKpUHKjYGmEU7bAGQLw9YgLa9IEDIhrmuH9/LblRG0guh
RNCuwKr38cM6ygl/9ZR8uyxzG2hu5C9ffZlNqFHAaAN2fNMUXDXAutzYBZDJdqRBHI8skh/Zc/Hs
m/tw/MKMMgIg63UryNM/cxIUBQPS2lzrmPgPwvmxZPhI4Bpq69FMwtAkI2l2TMmdWDig0gUhf05k
DYBI4pBRvBe3o1IzC+7jUZkqXScuDz9ApUvlNh6iaopGM4lDmw5eaM9WKAkLlDE+YJmAXxdfFzeH
/lp5w/Dxsoa0O0YWMANnMouo9fhmUOfcBs9LCf13JGagHZFnrvIa34mIkEikaloyTAicDxDEaEK0
yc6DznLAHlPigpblsIEr4ulyuoN2YcRggUu4zu9ITDLDJES5sdt0f7rFg2sWtzJeJnLOdoHo2zTw
V5WBBHjx/UVhBXFN0/HqVvJT2sWNkZi9FxcSsxe4xrH+JuLT14gqLB6FKkGTULcl447DTjxINbxJ
RYG0EoDKvKOaR028guzkGDdKMMpBApme0f5lZa7u0f3qZU3vTxcw7dxqo8+RGWe8aMm3UsKtG8Ki
WEuNeRsMQZ73uxLN4Pzgh/DdwhTZ43uwr2lv7483tosp5COLqGHCU5g8A6E9aKFq5NzGtkFkLYlI
amPDvkdZHXSrquXcaksWqCq367wAFvwF/0K3zc4ofDfy8ha5UGiXqTj4DEtYeEjQ6x93zRhq3nz6
04fZRo79O90jw8TBPuTsUpBtR7ieLXNJyFrwb3dIcxpSXs9jmf9mIgTB58QO/TK3XDKhreHIgv5l
JsjQVP4gfGh/hEtlUKWfQb3HhpjL6u6/OEeaW9r8DPQ3DEsQdQqT6LbPQeLlIXnujFS3Jk/2l3wr
hGx9HOr9igszrQ+oPV8z8bwiEfQSMYv2HffJjjHeLA67N9zFBS3w72KZQXOfVCVidjvpUOiOarR8
Q2FpBtIpfS4pELJhkS3vjgF0IICouJyGrN/I466Aa0397ErHWVOWgKLYK7LO0RooQa/Rr48yd8NU
hzLtNzHQ72On3mSfvA6l/4vRkoeAftsIaofgUFMfggsQ9Z0aFtW4bVyXga4RdTgb+X1nZ3EAahUz
Q+FMiktgVLtVaexPjFWAVarOa99KHHROeo15WEZ9CgLLMBATO6GsDsfUdF/E1vV6Q992qBj74XNb
I/L/ORwZM1W1jCzNzzpKjLE6Tt0x7Icg4lCcD6O8FBY4ST9jeheKZW40+Et3+TEGuLng5tr/CvMJ
LmCmvm+nndQjX8GkfNPLdwwzzL9VpEgqOtVlBx52NyTERUjizqrUnuwP5a8D58ve8WEtBKnSOXSy
2azMcrIdNmWbgnaniY5mEPIfJHZeZByJff5SDR6OUxOeTGs4/PS4IeUH1OUzhoTM5HPE5XOTF/s/
jScKUN0XyC1Hqs+E4ubdMu8zyPUJm1qfg2wACVHPGUlAh+lvg/hrmsiIEqWSsIu+AB6E7/RSm42D
S8/CGBhAGXIXWW3vKPbtPF/jNZ1Fi/SA6+SrsVQQDRYKfLpoPcS2wV1rJU9BtzxA7tG45KekIVc7
C5z7qlKwJELtf6OwbKNac4cGNX/X1TkUClpIsSXj4yIi2hKEl6GPYY9BKh7l6FbWf9F1rGW0r4Ac
xNlWbZwrnEFuH6W2dsuTrRlgPE/9tJojLHCBZk8H6X4uBEsXh/Pa6saqtoOxMXf1wZqXO4WHyUD6
DofNQtBtFMXu4x5Rf5q5HTSMzsI2sUPou08N53qPPSZVxnbvlGweIz1N0oAI2w+jZ4zzsuOR3Lbf
K+CaeJiXKTzSXaObz+kfhGbOzwmUVScnHo0j1nmjF1qTvfmIMA/0tJdhuQcPdlfqToFUtve2fUzd
nMdPpsecyyj7hANonBrnxU14Uadhj+SiWI9T1Gt77II8IVXKkjzUZJXWPcK5ek2HUn/NmbRt+ohw
FF/xxooufVjyo+EQGHRBA3UZ8gDuxh2SqWwgeW4A8TH/nVh33UlgbqfvfC98So2w3hhRRtR8Q40p
N6ytJIosLVWXwtke3e3SM+antbeyyZokr1fn76FWjsTBvUiFs/EzvvHufogG0S7fcSEwZ9WsbOGO
wMzZYwb1acrEH5JDzlgs30OcC5uK9DRAuS+psuOir4zb0QYDPqoe6zI1jL0wGqLP2wJfXdN14E4K
iaLAdEY9HSxnE+rK3a6Wkc0omhGjQXmrowWBx/Xr00+/57s3FkrCUSKyn/iGUy2x3I1pnIqosESN
jyc6MikIaHXA49qP6fdCkUxHwpDNq9Haog/FS8SFbUIjVef3WYdywmsxsmT98DfnHH5MGWlkDsSd
16ZotbbFweH4qORim4Yd6bCEvKUmFAcbSUodV4F9rHdfQi5sGcq3McfsZGAEbYypqKOYXt1wqOU4
33dmWrSh0qs1CBMaMxW94pE4fyiEOhbRcXSw7oymy/PJPPvKY1XWef7FgqWe8A6vC+BUSuGy/pan
C8fX9jnYXV2CVl65qzy5Q7omJzO5gmCh537LAoOByhs9mew1pHvmKZSu/dqbvm0nevuAMkm1M/Tz
4b9U
`protect end_protected
