`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
i6eAA1LFcgJu6f4SzGDuZnOjK2fZghCE3r+x25pIaltbxDMXuYq/3IBU+qlQS/F+qJy8BxJzXBiB
CKpebJeLHg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TeB0BxlTdHValqoNl6hJFDsH37SsY47V9OdEd6/co1d5lBXOpVa2PJ1L94D32BOlD6oStp7YtK/t
3UMuHzcL/Wgu9puPuqgXTqMezjUwsy6lWhoQBGbxX41FTDUh2YbsS5kTM0P5ll+wAjWzPxJU20pc
8Urw/r8vpnpMwRF7olk=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IrGqw1tmfeMBop812+Fkq4GjDBSd422DqHaz34Vq6cfFAGiEhAafCMS4jwcVFjRwgLIEh7SdfmAm
jFAQD8qLTel4BkfTr2onoEWOjTFtAAAkTLV/OBEGlRwMT5dILRH3/HtdV+w1hGw6s6hKDHP428BZ
DTsSGKFa3tsWnOjCykDob6SmkJH8geYjByy35+cCLgZUeC8nEpW7RG0EB4uff2N57I6xRXHeMFhK
vNACVL0gcMy2Y/baiYL5Kq80+klGNM2mhv7YFtvNjZxWkiFtd4TV/KnXadOwapY2vJtCTSdMJxvk
BcnWtlikpCXJGAh9nqnXwhiifnJiPY1SDLNnXA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Og7coOs4OHKsRHSO94YHpa3f65yc+oB6D8nBHGCWGWQXY9eZiCilGnXo89D0YXEMxFNCF7LtQ0O/
X47YnO4kaEULm4YN1dVlFGXDLGOt1iMeKzWgTyVBnDCjGOLmdHOJHY9DZoEmvvHWWVhIZCrfcSso
DAIy9csPriCNQFB62Gg=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ss9esp8vpYpUudYIe0XIcnXwju8Gr7Qnui//NGWfIPn3/6jkJaAV/d+8HG9TWbdcLdGV7qY7BlSj
9X1xEJ+kPI6crwt2WglgnV+g1JPpJPx2O1j4V5fTsuc3zo0m7+6IJeWAwHXBqGiDvAiuIAFRCICW
gtbZQVs7HHgidz1vIJDXEfHbGQLpjjQaqKmCSR4YJeFqIo9td6Zqa9wGplvY/S01PNUWdwEAIY7y
S4ZHwle8IthKhPoR6VYAzdt7QmoUVxnzTGRl1yTe4dxIy52k/7grM+gwVZhEIt9HUv7mHIUCvZTO
0ubyqMVxTu28EmvOZN5Bmlq9tj/7RtStvbX8oQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 8896)
`protect data_block
ne0TMjxIBcCahnbvK5x/YtxqEpiBM3HYVK5xhS7TqdEfNlbjGsQlSyCchaujlFELAJR0EjWImp1U
k2vjjJHZP9jqDucPo+zubpy6LQ/0deIihrXdK91VXAZ3qsLumIHoEhkCOsFhTB4zX9yE7HPxKe2d
LO6Ib8JiNtmxBFbUNjZbJu9mgIRXLa0uxclqfSb/fEmJDhs3FfU4WQpwXDKWyoTvoWQHXOFDABkk
VEQ+zlihfvNxQqbSLeIUPHEVKMmLvm0i1RxxN08z0Teuu9ys4PjtBiLPVYYN8u+nGaTDzP8oLvdv
p69LujK7RcTjVSLUnmPkTnyTe/Jvg8oY9GEyKeMN80irD3XvGZm4TsKtzj0RMxL1W6WcPj8bahnM
eh9195AoAFC203oo5hu63bRURxWRAyJZMU9YPKThBCOpZBFLDbrd5ZL2m4Ngd8uAVDbp47D1rZv1
YAEhpVCkgW3Ja7CmjBRrM2qZMvUFS85ZaCXP12b+Hhmt4UC8F3zGhGX47laJj5FDAqH1GbpZYLKU
1Fxpo2ztfPwYh8tsnTocfGdUgHj6sWouetPUJu5ZlJD5abHOCr0HlCALE+tqM9nS8Chk/cqTS2iq
0oyxLU+xzGQTiKaardrtcrYDs1iQXboVtpT9O5eD/yJSlFAr83NFRFMpnEER9qBQ9zEVWtSdPs12
VAKL3lpWKSua4RQWabGCmDQOJOW/QEn8zF0rNjwDuj4acP2dvy4xU2ln9eGaLF9MpC0hs1Ri8Myv
SBFeD+Pdt/jYBDGyaT1KTFxKX8edgOc4ZydYfd3Fjr038wm3UP4jxDIXcbrGiN4V+yLwBjx84YrC
D/CEidUrXtGBTAHQS+DWhcwCbr5wGoQHHOYCsy1tIfY5M2j20PvAggiFgJlsmo6Rdv3vMLCTttin
mI39HT8dJ6nef87ZQvoGVPYedizk5c9YWmiUn3e1e8br3F4z8uvMd6AJFK0KsPonXYG6s7qCoE6f
D7R1li5JkNkrkhQDQJX8Gxl4chQrkL42/d1chYmvmLKX2Wn9lMXXWzmF4Vn4WN7rv4UIdN+kyXCn
cRfNOV331fimAkbsA5Dca4Nmh9ZNUxK7G2D9nP3cuxEQi7SpNNg3EfPUYku7yshuIRwBMmjG+dBK
Ul3OazDPid6zKiHYOQbfQngd3mCXEIz9izQx4Yiv1EkT8/udadWjZFBbHc1GwNrowF6lRhY6jn4n
gPaW7xey3tGG/duwwrlAayJlNZdvQTbJ/xZdnCM+owjh3tFba3i6m6fZkv+wgpzZFeT5OTpcaazA
Oef9J+KyPUNEBb3kUSqJ1v3l4d8OE9mwuPQxZbbg1g6V1Ji6FQ+qBYD+a7cIKA2cspRXq6HcRB78
e5xfjCIaYvp8NVVbQhoiYBjJs0I/fnw9Bh0UTAVoXmj1s9AJpJfjGzdCf+LSypVNJvKhjxvqIJBU
jKkaN3p9eCZBxhYPI/NEOXwg5XLzqJeLSTYnkPUuFqtKnEfIS8rXwaGnI7jq9cjdUVFjGCaYw05k
uqlPQTgQ/Hh9Ct4HxQqQJ8ypyUj8daHp78Sds0kaLO4SsVCu3inviq1eN3JqSryUQtJyF9idnKL7
9FpN5m2FJOas4/2l72g21JU3lH6wdukL7Ou+Mh6GEs8UFvdiUmC3TkNU0OKLaUQ8FtfDiQp8jUow
GnyM5fb32jbTnMqqbD+DNI9oBDJhSoV7zk9tezSf91D2db1yCpohCeHuJXb2XdgUJkUQjARp0+gj
CVVjBdYdO+mTnXzv8oBP4e8Ie5l5hO5IFZIw468IiVDJfPLTYCt402KNP4XkTm+pmBM2nvWPowcH
E+8Ix9/blagg2A/FyZ6z3uhQV7Iwz7zWCmiMxgtoDcGRT/P5n1Di/nI8x8wXV88gJj8sG1/Oz0jb
SBa/m/967yGTCaMnQTeZSL5TY8mNRPOwiXWgprWneaAsFI2L7Sb8W7BBJrgrLgX/fEoEjqCdt8KH
8xaVfF6tChk1nFtf+2KKAQxKqi/LzNMk5YJdhRZmb0EzWhCtnOseHspx/nIWm3l22GKqicu4LKxm
I3851tFZkRGOZ9FtUAr5w6ySuBzYJReaOmG+xZiy5DyEPGb7ZPcRbZFLXdbI7r4wTUUgXcTff0pJ
+xV2hyvopPfNFKZ4GCFaIIrtHy+YAt4q36ZiOFwhdOtLu6yLS+z+aDxCe7TwU0PpN698rNnqqZkX
la++PFlC5yUbO5jfSIM0jTpI1sKQ2t+pY+Ues77MmJhyw2nXUGyJ1TRa0Wv8tFVJP6skDDuDqItK
XZEzqeAwID/40n5r0TEBOsVVAvj4q5jA8HYAkWculLgQ1LyS52BjrQkO2pUng1hpgdCoI1M67if6
zAa+vSAOEGixpze0rtGBZWIQBtF+t92b4lo8pHLAHIc0E26xRv9EcICzyS8Sm0HwDqO36aQ1hYdg
JmWpz6L17qlwWDmEilkcU84lD4B3rTeiv8NM3xNM0LsHl9qMWXWAVqV1QlQOBEgTxAGb9RdA/tge
C/ZT23Bi6n6NAgEOklAkuu5LHATmJpDdimrXh6bLnZBxRuRRbA/aZBB6IpiOWoXZQReCqAHpxRCS
sbVPK1ARDUAi5hX3DTww5LPHw1Q0A5jiBVJi8vN8c+bIO06J7HMWP+j6mgMrGbD9GFk9Ri2I43Vt
vldsN4G0RDcZwBzCmiyhsCprEWmQxgSESrRHigZC4fK1rQH9z4zI2AzQIUHS1y1QfQ66FBUC5H6X
yy8rtEBuQL+4y+BsjBsZtF4pUKEeY6XbYLV1K6Sd69MexpBgoHtLadH2x2wIhj1HHZkwpZ6JKlk4
to09bIpeMCKkE8g4tm/wrweFkm+plsxbgJmKtX9Q/Y5veVI18XcXLXylwdquA7o0aE8bm9ZLxlrt
4bHfDocTMdYXHhHeJDTMC3iM1yYN9LcBAKN6RDUun8dwuqIa+Y+DTJ9XbqjRDqBzLOZGtu86aiCs
VSwKdxTBddcxIIORwVWu/8jluQMw1HBCiL/kFQcdnT9yvcFFj6oHj6vRUzmoC+ct7IPfejgMSzfm
q0lJvH9YI9/cJF5cRklPlLSYbq2Wj2zHcGZk+not0cEpOH8/b9P4gGVOLawz/RtK6+ckyydTdDab
yDbtbd24ILA3IDtoqhxW8IqxQRJMTMJjQXSww11eNQmk8e1M/nsvye4NVbzwhwE0EcvWUAC/y6Rt
LPiBQVY5jX4mcGW60rSoMgu5SXZptql13d5nsDtOmOJFiJrOlIuGrso9f4Q9GXRJUf02yJP1jOxn
x7KdemcMGRwMD9vLRtuP95PB1P7ecVJDk1gBkl8vI2GPfGWzWlxWWZjKy69XdYQo1kY8Ln/rV+65
yj698t9MJhIp8rLHmhl6Euf66Bcu0fKMhgw6++uDPnhYH4qqjCJUNSFtGvfuzfcV8YVYAi4DfjCy
oPtnrmD3gFb36J4v0eFNFgRYXkfBxONqAsnQAw0WycfbzbEudMh9P1SmjiaN/E72S/qqBoYUSucN
XBtzoDznNiN/yG/PS8DOCKiK8VpfYGMlWyV0jx/AhZh135ireX41StU+YvvgOaArDAyNnqT83ohH
WT8jOrsvBHftOrVZW1mjA5itlCso+L0kGI0cWf/p4ZHHaHW4HUJx6ha8ZWAvkDS2Z0EzM1ARY2mU
B+GgVoh6FL6VuPCBPqGFA67P29C/yKnNv+7FxTFUXPAdEyceASTBhQsNFYwJghP7Izg4FMDo3YB7
AJRT1bbtZmitYrYHUeMXhDJ4TsujJlDJWED26UPGzvK6XLUKgoeTE2b+etg2Rkao0Xn0Q92M6fk0
8eJrVJbdhNI+4EEtRwaBwUKGDksZDPCdC/DU+QpgRWapW2LVg3zSb1fs+1mqR9IQoUseBDx43xrF
A4tPcQSwfx40A/NaPG9080/n+DLlTUrHc/UxwzaFVKy4IRPIHAgv9Jd253gJE/jzqv+YyM2f2bgl
uzjqlYjSEd+fUrsV8BmzhNqAxIpbg6h99gVSVb/N52hM0gXJy+Ig2poYXXrGRSnRsl7V5jUg+C5u
IudzR7whiaFlb5CaphtbqPLFf7ILGu43Zh6BllBxmD1tZ9//a8aiBsg5hap/mpNFTDWxY87ljxpN
ly7PnzNnhiiuFOcV+SPsQ06p2YMmxQXecQQq9C7qw5IaBred0772PUcnPoX5areAj1k7bEwpW0ZK
8SnLPcdGUMpIFJXB+NhrmWB2ZK7Xfkv+0UldaXuoT8aqYwAF4eUienT+zIYxPk5UyBIbzd1XWS7M
chcBi+g1YTFdadvGE88uCY6xepzjf8bNzSr5iOZlvGArVRgFyqfbQ8NEoBHJ7VPv4aOYCJp6ic1i
u58GPNxVLaySI43C3im+XD///qPSX6Ql+CNpUe2HqyVfcdkh+0l8ivHFlj2DXuYYsTdF/CBP67vb
sKwsKyIwlVH5SCyDWnCQONAwwokNRDfYJiMZsspcjcuPWlCOxls54jq7F33Sc5Yek9MNCSVvnt3T
KCpxFOR74zC7HMPA/5mUNRwg7gG0w4hnIcmTxKEb6DYssiSKr09R9Td9rwW1Eeih+8ch2K6vqHvS
/7uTlCK2qlYQKE4sO7MAYUyaG3WIpwcR0OQm6LdVpWipQAeRD9MAAup4dCRD5g5sje0fY4bHlQZZ
emIZiHLmjF8w6cbYoIwABnBxf2RoYNjey9tZQluJZfCRebTjGiWif6y6amLWRXv75Tl24WqgcgZt
F+23OxfNlUEfsTijD2vKJBjpo9+tYC6T8CDHX8ztfEiM+wJ6mGwZfHd3+dDJwiSx9jy+x8WQlpVE
541Q1VJLpDkZp0oq5zoah1rb+yxEuKgZU10JggqrQLAWPvEDTlwPp8AMGrsAToors+c5itRAAA+z
VEyQc8bJisAA6yQa9jEtMGU/HhUbHLcESYerSEtNh4RiddhAid9kOHTNdON2lJ6VmGVbXaJtF771
8H2bUcxHMEy2CO4lasuPfbkHLE2EWCA3Q2lFNdln+DWaGcB1e4VTL38I/HacAPK3YEWWnZdu0tDi
FkB8nweY3FK6jwcvGb1yY2nTQu6Pn0UG62pDg0gQq58wGAjyke5Oshx+uvIcM3aAmB0L5DdyXmwD
gK0LqRH6AyCdshwj2QwN29fwb6kCfrKdRnLlVfAfCIGbDJtkWwA+n/6RwpPgcUPfFoAn65rXBGgv
xXBYL9yMFa/Zt0B0JgncIKfvkb2Fi4eu48piniqjZsf0g+uoTSZ16n7K1r46f/u/DZ8X5iRoWTrm
clwZzyBjo4qhydm7GdQ+cahLVIrVtSqhEY7g2TfBzvAb2PI9FGmB7Fe0MWI1RzeMyPjSz512Lue6
MEO6NRPhtYAHBOjAJqBnwL36KdATymZKBlbZ41744GXwMGcqWY5LVsHDYj51kchFDHms2C1IwYB6
6lIeeTQKGBIOecs3pwOTgf49rkOX6U/fad+5gfK8EjuATPB4XPD5kVDQ/z7vFfE3Qbhc7j1QKian
zQRm16HJ2TyfhP51g78gyXqDYAnATKtHoy8y0XkhII2dvlfF4jtC/uLYpOcnh1kderGDKrPyeYfe
6ctCTuKWIH133XY1E01mt6+vtRlW/pYJpVc/RADbFYaT/TFKHcmZbfhVHYwJyguSZ9VSFpeE41nR
6jHn6TVhr99FhOHkz5DmDe190xckvmKYPkM/+qlEsMXKA/i7zF2iz7KyKmXVYKwg/NL2xJBV6qLy
tgmL58YvI1nirwh4K8QUIJ6VTUepFbLJV7TPKGQ7lYWGUkPnYErvhT3CDyiBflJFSWGZHFFk7GbT
u9WsuxGwQ64Is62k1fOg8DWtLSN9EG07ije1WuGbTzX/arbk8x3cdHbsuFzy9aYTesSt4OVfs72x
IkK4n+LBGxAAXW1cvMSoMs70PCNY3nod0D90GkY0YRfyvQAioNz7A2d+LP6bWfYFIwhIuHvL/efx
HSEfg8pRb57GJe9oDBZ2Z7+LnwQ2+Zfgyvz8dTNYAo3NR4bcJxBJcJMrzkQJwF55rkprll/udgm9
/PQD65IIuiEX1AUpAs91gVM3H9wvalOqHejCWyShRkRo7xFQUA4tk6596hCJ0KwBIbIRFVSlDj5j
RJ9nva1mgT2UujubCW1d85/NIacUxe1SddOdueDFtxtoAoidW7remb+IbaQB/xiH0wHGz+2CBZC3
55fR51uSQnvo5tLlQ6vDpExMM10qHwIohEfpx346TEMHC3EmfTRrUhy9jQo4fBfXRZyqDxwpIhQX
iWPx7//GQipb1IjA/RIn8jnMkrf1LFmDEHG/V0JVxrvKoMlGSIDaFdEHC5yJ6RS7EB9gTxWg/pp6
XEDVYa/gnfS25Cn1pklgEbgIhftWc/808c757zMxzyeLufH9xzZpIsjrzRxGU4iqO7RWJaoAkwVk
NNhtoM16wk3LorQ4d4d6WXJ9GbdZT+vURYDIOntMP/nMc12mISZWac+9AAO/bZOKsKXeG0jTfbaz
1EJbqQ19M8FXJo0LW9KsXcB8HnrpGjdQQWSK2u0V8AOvfWsJH0Pr4D5fbmJx5hXVsHBCr5e7dl5q
iGzWWt2vy2XDhv1D3hEnAgYI6hP6d/fpnU3Y0H+UTnlXbSlVsiiYUMp8d7i6GVnfmCo8zppQP/iK
Ojtr79Y6dbtc8jgUAjBVEg1TqctHJwJzCqntR7cNRyodwoSJhJtRUykVCgtO5fVGIyrofVL+8h5u
TP5wAygKXLQLUDhL+Flzt14bw4r3o+w4xrQw6zZPk+CC2/7saJasg97LNuTZ3lB20OW6MMoBlmRR
9VNsiaSfFYJBcySRND8OLPZH8kiXs2FQmzhuljsb21cgcZPvIWit9zDAeBNoY9zafFW4K/V65gvu
jHWrgmoImNk8kM7c5d2clKD86ueQSC4S1xygbBsDtuecpIUplYMjZNnJAOTAyxaFU99BmUXhmYwk
LV3y51sZUz1gx8IR2n0QiEuILd7ohHsqBqkA+LO89yiDmKS4Z6rE1wxkUcspaLqe872If4vq6x65
Dw+m56AMsX/KutPSNC2mPAT8UgETm8ujBroDsEqqieh1UchNlMe6SwDWWxvhBZnP0FkNmgjBVYTh
SbnfhTNATF/f3I5Nmg5AgzwBOhX8gPvjzKvdOopEPnEAYpcM1jevPBV31KteWhO7Vg0YfIAafoDg
L9eQGtDe/ZBsk2RGij7Yp+8V8lUenueFi17eSILG98taRo6QCXLDNK8/Q4wCA5kx4HUrRyFnyOPc
CgTndxKTccBSL6BNMfANR4xFzpD5DR+MU9CcNa+7qT28XKj+yGJqxMlQ1Z5vvKV/gZ44xKjSQe1l
7l94uhCrRvyoFj/mIGq6vTSXfZl58DW7EJOPQbtW3WcpyOihIBUB5KiwIe4xMH/AnO2MpV+HdcHR
JwB0CeiPbJjgSb/RsFYfWtuRSiDd6CkwJ/nPaFN+ul+kL5COkWpT/qcL5M7sse7DihKnrPvyEAWd
wsREo2GxpZEnCL/iJA4dfRJSsUJSE+rCjSOl93k5iIBaX8hpGEO4ndgZgLHw4iH3YT7otGQj4fH7
sKHpJcSVauLT31s53kOuD2cyn8l3wn6ie0hHNmKZbqvGW4C4I7YnPliUzYLZoVza/6wKIPA7ACy8
M5bfgr6QiHLc9UuVAJKO7m1+7Gwl3EKPCU36B+6pKCG+QQu34MQuuYu7pa7cYaggvz5EWcaFeVB2
o6i5UYywm8luGyYIJit2Ic/5V6K/Rb8W1L/OF6DnDTFSfP8vVsBnrDSP4L0ISgLeXo2z9FfWz+BB
kotaRBBU6LcSv/y4Jqvq8zKVtrRiasf6ocRwdsyIOk/WLj4e5STj+wKIJeOKBmK45GVVm5umgp95
VvX+3yitweGmocBdarxlf8p1qt082iCthWqe5mDOTrqPbA3IkGS001qVLT77VGOQFeyn1861DbVV
T1XTKVWYKQyt4DIUN304WGRHwU73YU6xm5AbQ18MFVvlPuDPLVwmCgJ1Q6TY56Rj8SIYCjr/LlnO
qQ+sr/AkP0cebSosxaJgJJPFulV8YgOuJ/GkMvNX0H1ZRf3JOJgI6lHaxh4o/NScKiaB5v10oJPy
DmHitFOVhCdbYY9ysssJDRx109uVdNLUgPTtKPwDWTwtl6IAW2PZbfxFixLo7nDqRrdg4MMFYvUD
yj3lsRbNzZZiJAiYT73wqJPALiNuBAfx3EbmxhfLTT9rvP8cbVHhD2fNJ2eEq+A5KN22LjsmpRY5
NzbAurUbS3BT75lnTN3vo6z+gOdBYyhPWZq0TXyunbXbAD5asbm6zQREu2mWWuB5uPG3XgXwV2T5
z8b+rxK+EnXugYkBFlvcOSNh1+O90ZqBL5D6R7AtEYp5Iav90YU+cEeST0GYN24+5aoItSDw2XTw
5aBItdzLujcUVKD2NkY6Es3Vpe1NqgldV4y+vGPLk6Jq7Cl5OHObszhsC+ub+hmYqPMS3PHK5x9p
HVgSVpskuzQfVOYrvZIYy/DR6C2EVjIMegaLHuUJh9OeG5y+6fHX754OdPrlp6suxISrm3lqrFPY
WLJZ1SSHK6ESb9TyM/BVan8U9t4bm3k4KlVGn543I8Z271VgrKTXEXyslbz9LpUTrCMrGaDOCLxd
QcDGFp0YeZZgGe40F/Q0kLs8DhAphm06gNgingijdexXxGySnUVMN7eWFMXhLrgi7AqGP4QQ9ASI
wxH/911LcjbMZGpZ3dJ71owE9hcfJCzWDcLVorT8z/Kzy1IRg9OUaTtIoICdf1DXYCSgtOPPuu08
+sGr0D5/BFHuKIedOgMY6aWKOHsfugF2L25tulVZ732wFzvPkOC3gMh5s1g3X5mklfnsp2FTc4ms
f1W+S0VeExv2uBx3dqra0j/FdKiWieFlfQz3ESMEttra7LsB6qN6YWA6YPHNZPbReqe827iZ+2Zp
5jTAz7K2wE/ixBUE/YN0nFAWi7VYpPi2d8ghBqX7mMYrMO2/xepmQHB0coNHlT8L6in4FRlnYmNk
PnPf1ScDOvGgvWlO9KRJGAlOo6s2/YNxGd/QHUc5bOuMRqNMNePyeHvsce6XRDPwCe53V93kpnZN
IpnlbvfW58E2KlPeYdZdzA5+1TEhkHaSwtwTHKGfnBdnay+UMeK2qzFTK7yrNm7XZpLDYLBtLwoh
IrTIQgODsiI4aQ0X57nndaPOqTcrVaGXoxHgmnuNBmadIkijIaxcvk3TZuKABKTDgtG6+nrD8eSI
W/sgMv8bUMUslcTZNauQRT0Wzs5/p+qC0SXy+/h42Yj6BHQI3Xue51TtMW8CskbtJtqr8ONETVxr
xgkPlgdwNE3B32zUW9TrKZtdJEBj34Kx2grYWzvy7gr1accJxnmX/qX0ZG2sneY+7IqiaZxpj5Dz
MJW0x9789BiLOaWWB1W6lK2LDCHOvXzplj0m2aASyxlyDXzccOra7ROYXw+bWDm8CPk+wl9+C/TT
Axu5HBn2fVckyi3onv5YVIEmI7j+o4/t/7zY6CR/Qoik9uVbqgNQhE0p80wfj96OjdyqFiZjULs0
H5WhseT6TCOIeDz3tf7uh8P2q1OAlaNLXiagU67gwB8FcT1KSbZqb2Mw1u+tyibq2G1ajXus6FCT
nItfdvCU//yICZ5Ogis2j+mmjDBrbUGOdDrjx+8clvhu4kcVh+OOTOJUVCyRRWTNtASJ0af31pFV
3StB7P0O6TJEHWWr/v8XuqmlZhzae/45qzPt2yudz7HqC8/xF/nNPA0BowQRk613xnatsexEigDK
1yrcBpGiMz0mDujnqzo/y9WGtlMRhOhIJQtMquEt72gLe3y4czu1vJLIo2UVhs0xHJKrm8ATmzkj
y4G6bvLfNAbMqt3Wun+mjT3lUPz1ByDOF8Fpd4ABME86Qsu9qS+gCKWhQLGlW+d2WYkZqeM4n8CL
wroH9wOoQiuHJWoKkzzx/I6rw8MF6/uCAfppXqLLYtpJCyDajgomtNwt6IxOTVssW+8zW2a0o6q9
c29ViCMpwbkFAkjRU8kWDer40xOx5o3Obp2h/ZlvSg6PdnuByZgqAhF+u+v816JmvO6E8povkj9l
XP07uMVRIQ0t2wLBFB0j1mIpWN6eYGymiui8QP3OCtNgtO9+vliT98yN+YjF/HzG5sKeuMcbwysr
BgFHUa7u4V82rRyYTxQYhkSeow6jUqwZRH5nzrrf+iywF996KXE3hfvs64h2WXvABoRwbxvku2qz
jIohYjqQmXXTf0rLK4MrxMNh1SbHfVCplcf1atZHotzRAGXvXvBSf78Zh+UxK8cCi4ztC5Oa4s1V
aG88WlXb3tNSzIiZcBFEj3VBumyx9xrHqJN5x85uQ0kvgqjjbEQdtEqkYzF4l4lyy+zWYGcBD5Vz
X9TuST6WT1zLRV9YqPNGoMP02fh+qXa2232fCT3NP3SJhIEKO8PHNLwk45Ti+PM5xWq95LadWx8x
/7yF5xmb/kwYIebK2USsAcqWOH0z+0XA71NmIvyarbB9FVg0HN8qjmJajjZG1BrkRFYmec035TmA
XO9vtI7xqKVeo4/g/gSCVYxDTOxKCmLNHlTrFiJYvOWwh+SdgUa5VmCVjalIk/a2Hj+N4N1yO1Ub
vhTFt2KHnAPiR7NeQumpi1gy5YujZMt0Gk+GdXwsKkQ/e1f+GsR46YeUUi4b4ldZ//iG6uaYTlFQ
SHj9XlEhfsUniX21b5mMfxRCluPZEyZ5wYXrpFqHyAOVVu5RqgsOpMu00JoONBRTuATfXrOpfgSn
WfMVKOkjtJkVMks9bc7/A+qDxwfgKpPx+1e4v90ns91L4U/7M3USyg50NChMbKPO96PjbeuAYmSx
ezpB1xzzKRLrRbGB6ebHuTLCEqlP5lmH/RZWhpGsfyky4L/day/6f3FRkOG9cGUyp98FkBdYSMfc
6zsc6UdG+uqHHtlJDpE3C6BALtn+cynqOsIm+03F44/lupqmR5fSgOfSWbyTp0LPg3ZvnwEJ/Uc6
BlhS3Jxb7LwukwFIM0dCrwuaFbLl6p0K/bsUOLhLeF5GW9uKSILiJHSdf43jtQUCto9MujKwzhcZ
Wr8+dk5WP3MdELuFxz1/vtBfsncJ0iFeCO/uLofhi6m6ff/y10LjhAnnihMvCvDfE7tpxHuXtrQT
AdkdjObuSsbUMDaaQXpodlnzRs4S4iFDfBFImXcV93Ssx8xzV4I53la7s7ao8PbDSQI7w1Li8Vt1
WoD24/7m3TuYHNjqXjdRJ8HZ+3ft1L+t4kguEwm0/5fT2GzOxUXpF/dUkArFYOmxnGrefUY0MUTX
F8GKpDjZthsbXs3SmFoM9qcnDeMDJmDS+0qRy8bkYPtzhDJXAOYVDlHDpnW2r183oHnoRa4WH5oj
YesKiGE/M8PAQfCDKktwTyou0/8D55n0j4RkSzJZg5JlcZWBeN9b5VKXOyD2TTAFAD8k82TARVsK
P7ifvt5Q3BFGSA/7L/FUlgRNXrdP2MOYwV/XLswz9iDYMXBSUzUeZZ3PO9l6gpFhSUwNs3BG0f1v
U9pVUmLT6jZwX/NNeYH/GDYxwekzFJMOshxCqHAtC7N61R2jkvKqxzJZ5OucNIHA0vizU6aswSn6
i2+JdBqOMLGuS05SjdqZJBgZz7n1DhaLrSfeRMsV7fykq1BdSEsjUkS6J49zrp2R58lXuUOJKqAn
FBb7Cma/ccWKMnEbU6orj+P+M44Krh3JsdD+ugG+WTCKWf9lroZsRjk0A/WMFQODXbbmoT4ALD1X
ySJ/sj26AQuEpE5pVzm0YDsWNqm2rVTs/GdDU69VbsMe+qfQvL6z0gUCTSXsgDxVm8PiXpUxsItc
P22R8nKP0hfEB/B8kZ4PqUO2dULjkQGvfYdBRoY2kcNpYsCMs7uHku/YWbQPbDn6R3qX0LsaKTls
VskHEQ==
`protect end_protected
