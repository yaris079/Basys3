`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
c1TTHaZmax2QKFmq6ZfGAAFNEZr5D7u9LYfN2IPUBN2bR6bIexzmtaMe6ju6bQNChnvkuKEBvsrC
JnyvdCEO5Q==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lJRk1/x97X7IepQXoIghPrc6o9ceeaKrWnFpDh/QCCMbb7UmZdL99wJQmz1/wqn4muufzc6mpKvR
/xNyiDKxDogJH5i7G3qTXasK2lwtde09Iwb8aSMAqJRg4SAiQhjtbh6eJ3qpyrKcIoupGdWJN7yr
HaMbFZ7cWQ5Zqfd+tGM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d8AHdSrf3OlgkCD7AoZq5M4akFG+uETRsV/gpODbalJSbRPa7BlKAd/2+3EY/PdK4yH6M63NYsJL
4nRAFpA/DIQEVsKpdTg8fDgJWc/lp6xF7yMSBOPwiA+suBYyTXCPnDF9/SFklNg8hloPLXnJxKdu
K8ooYPmvtKuJXd6a2OxuC13HzQ6chEqyDwOU7iF4AT5v/HJI3V1t35lJZj1JT+cPZscZV2eBuF9i
Pvyrni43zOrS2WzS3P/tmCCD76IxCoMWYcjY6vqVJnGZG4Ezr+Bhj/wSrpU1Vs2vV8bCzkuY6OeG
QbO7ow7OiAZwLcJ4YH/2J4p0UODAjEi70DNfEg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zq5MPi4olNCCndUD4dIUdwk3zjFELpyw6CFULLJjOrNUa1nbBCm1u7tXH6nfWZoM/9a+TgBkmCYF
IE6pw6oM+tpQAzrpFyPm7uQhCS2F3HGXvSUqb791MKgNCm+kYtx1K66aKl7GwgGaOLah5XAtyW23
0P289DMGmg0kyUGRbp0=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BYtlVg/S5cCZse3tcjyy4jEC96jcRjBxyqyDAD27MBtj0oMEHzg2skabd2HoXr9URYHf847fkD7N
cnKEkoHsNYhmLsjdMKjMksWqzb+BlP1tA7hMhaXUyIC/LMWLLBp1A5ojKicADs5p1KA22sFB5NH+
2YBt6xtpq3dkFQ5DERNomGVpgduoilCTDaCBqAdgjVawv68Z1dpdowG9fV9Bz26O8uNqI0ziUcXV
7c3HuzcH8JOECtBDEjaYrwmy5nS8ycYjhqvppUftr34NH5nV5y5kz17EDx6lSsdtjkScUEC4vkDT
NkMSV16TEWXoJ2INxR4IqQU9+o2nP13scESCzA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20944)
`protect data_block
z1J7tHBefdtGJk77LEvOxW3Koruv64pWSo+4BIrN7ZEiXCKdki0XDZbTPoNgk8h2bzP8FXBjv7IH
/ArjS+1m1UL5rM+gmw/4cnNsUsb3UMUfu0QFuTAaUd7EZVuE+EBi2U82FV7nOS3ibaGZ/oW6tTSQ
QzrHMMiGIVO0+Mh3NykaBKRoSs2NczQkmJYxizaWHjhQuJ3nz3sSr26F4Syyhc1b2t0FMfsB0Zmz
VLR/Zp8XREjtJawypA7lgNepd3GcfkrhJvxjUPuzzExWHTJ6BrITYBEtZRyuTdakC/+VfuNCFeWk
WzzC2L4AC2D6EFUM7JW/uy9TyM1XyJRyPa0wYee8ndsrBrBmyJ9xDJYNKG4ZNXYrAqH6MGaYSVWr
If/+/P9PIM7EHr4EgwCuDa3N+sJBEteQDnOX9fzS1+5kYT2auT8fvN/6jgbjCGBMx8XAyX5kd8HE
keycPgvMkZ1R1J+D9dckAwAVEASz/ljsG3XXWn/eFmYkyTs27ewtxMUCDQdn/NEZDWR4A+t8FfmN
H/hTdXjRFTnqKiw/tCV8zAhnCqCDbwe9a0qkRaMCdhqiFiS4D+C38SCa/WbSAWajF+wXA9VFkchf
l4RdrQygtxtpJqp24ICVE9zZlluvt+SSA/OlE9ZsEG6tYyU+SLCDvUhEGu9pRrE0bw4Je9IJl/bx
o6o57lJdZyqcNdh3xRD4VeusfGPzrKs0O2VVjAt9elm1nt6QpE5MbtTtQx/PXrDNdt7qr3aTgmfT
TRoWWIeFHMvviXzzBAdUCUO1sDgUmolw4vVo4KSuMba0xN7OSHKjxmr2/Ns27Jh3c9ehu9wv3Jd0
i2GMG395RbBG8M/mfh7ksSMMIJ+M1juhCZRjBUqFGRCJjzSjbXebQayidM/QvFqDNWaQgLWBpvxK
t5V7JglBKjbmChYQDSZesmmZ/wtpoJs4F+bPPFDRiJKpDN32O4lLDNzO9JS7DWZ0zitTd5YGFRe7
QMob2HbzVJIH9Sy1mRILAfBikPkpz9c//IRZqbuZOz6hZpqFPDVkHFRNuRHbvCuTuVa9gNbav36J
EZJmfCuH2fo3IChZnyMGKjQdey0oUpOzCUM1j/5Trlj7u1Yc6LQS+TzSSNam/E5OaOunODzWOLD+
UaSBQ85G6pIO0KksKEWTxW8TKGv4YEnU6HSKbORlA4suyXLFW0mny2BSKyZ14+pYMoGz6ZWwD+0Z
CXRLRS23P1taP6U8C6fpkVzcd+Jcc59z/dEf8AQxgVzRP47XeL1FyZQXHHFRJi9KNbRsB+4Oc+Xh
3a3V8yG2SfBGZ9Jz/tQrF+HO1BWZs81XN/w+LDdYxAsZPoHvoSoJvhhAnxnCcPDIbHzx6vnN5/nT
JYKg0h6THwMnjeK7Zno96X0qiSCHnRBLyxAbydyj4BUPSWgEBHEABRzMwVRtEkh+1q9DHVlbit80
t6ikrNix/Ocn3MK1YAwp0jVjgQc4/V1zlU4zbBPt5K65obxCwGNJR4gHqmKz0z8/fmp0qwlzqSFB
LiFUFaU27wYjWI7PWp97BW8zZIUYfJt6U4Y1IQL0y4r2myw7wRZdRCho6ssbjeiw7V5qMUaOcOFQ
F0r7j7000kIokqHkjKgmIFY3XFX4juI5o/wtFS5DYj7/knYFBRR2eHNf64qUjCqmsPfTht/a9MB8
7rgPNR+04WUcSsyrncD/4eUiwtPJnUwMBNXqAYO7P/oospZemlAbd0UJmE07xggD45137yewOB/k
Vx9v1hiJD6jOXV91pMGdFekpiEC+d8bFmkVYjifQvEYSBUNcSrzDFEargnbBvLfnVU3cJP90rWL3
WQB+830JV3RDKafZYCncRBbjMTgZvz04RI0+ONqScfd8LTIm84HKKH+crW1Dc+iXhYcVwqEGLr55
tuZzsF3J8o2M1wt0mTS3vEEbZx0iCcaOIuTeSHDTaIJBnM07IGxWPzH2d3EPN09Ox/pq6UfXlASn
YjcBPkc3CN5yyS7xKJpVZlvp6k6I8Nu7AIIVKLvgZoWNIBnfnn6OJLh/VY9618T0SorEEHB1bTkJ
hC+hEwqUCJzWU06NCXAFCUPjuDrgQxCNbI5pf624D4iNl8VIbJFRxiE2r1/h35NOZVrqa5UZo1f+
uooo5R8A3X8kNdQ4uDwcdNCl2TtxOw+5XsT4skmqsg1KFq35KE5sWsC6A1Cayb0vIm67F3WQaQjB
yDgDPHk34vZR/Ak0o3y7uct0KJLHwT1TFIC6o32q/K1/j/aQa6/qZotUN94YRJl1gu27w1fHWBQV
Yb4QiYP+IZ6t+FmUFeTnFGtS+rgUz/gZuYokuB4Z2+ZvCdncX0qjbCw2kRUNJ9FJ7mOg2OcA8Sxi
uPMB7+PvCFhBzmiKYsjUjBuOHDZt8yK1+zHIg8PiGIdbVgwXkAjFy82VmDhEVSvrO2d3HCqHnARX
ZXwvBm/Q9QJ/9KFhtUNl8+fSIKmi6Jor8Xu4y+C5tZXI/CbTUapKTRNlvcv9jHZbzjGqsL2ys+M+
JNMDLo0q4AwWvPfyXw6bFDfvcLwPSac7ac8eMGOd41a0v7/GJ2gvTG2d1UypjXfr9n7jIz2RMHqb
kO9LsbszqRb6OWwBVk57M2Ou/9VMFIOXFEEzKVw94fB1Hu9AmIqNkjaqZE4wW4P8PGxa+EX8V0oj
K/y+uUmAC/jdytTSpLMt1iNnF1nNk39/X1P+X0mMhVaV8JB7H+7/T74tzDMVCD0Hb2iUW1IhaaDs
93XSZWfVl4ihfoHhsOH+2bzBcCUBU6VIOb4KqyEL74A2aBSQuDjz3IUgXiTTTQWGW5r1I5ZZ78Hy
EM+RraOms4LuFlc2HspHktRaME/ktyDcfM63cmwRJ8EGlGps2N4jbFZXu+LwTtq5F82vkt5PLb8s
mdPXS4jFIo1jeo7FKvs1OnzIR6Kx+c5Omm7qikbuGMmcanE/998yD9rjlpl/lRIPk17vqXO4hwpy
QdJOVEJROP+uA0qgtk1hiodKGIhsJOsj/hO/8osR8rr6jGCCSB/8bc21Oh+xW/aQ5D3YKhlrPKZL
x72ykkOJebZ6k0fG/EBnoeEPXtIAL21OuUTMT0/tfcpyy+4rFJXSrnqenTjaFAIPNztBFoi/AXBo
f+BQgtxigyS7pGAVoOxupTECjrzlNfgWx5/9P2bzbSLMbF3e2Q6qYc+PuKnd5j16G3X5Hsk2CBgT
Z+3shcIqtZEQszrv8nx5vV01DZcA1KqoDNzSafVqM7nw1N4N5uvRvLRaIG2is3SpfKwf9ux/oRD9
BMNjdB0LzeqXLe++UaxYND/0dW2rPC8OCLVCxFVfv48OTlKoSKRIMxbpEMjXUoluqZYgYloO/Mlt
HXxCgzZ+W0rR/T27jyMY2dDBN9e1hDHxPvD/ib1jfJ2XcOUvWESfOOYPMThHVwd6a/DoJe43c2v7
J0yGOTeGSELrVuTX6uqN/uH24RsRw93dUB//FqaJqos8OYj71vyegonH83fdnzt7MkhlzudYQJDm
mqihgVGAY+hX2fj+dKIuEbrCpB0SpiU1WE5jKu+Y/G6aUxHSX6zDnFuF5DRd9O0YFAaw0QkAfBon
CzzQ7gOQbbP6LxroupoK+K/fpWKR6qSTHvtSk3WJSll78BIPE9vpvdDTAiEo76z+gkerw9ARYzXG
aCVOtRK9FTkBalYiJYlLy5h9Rt/yGrDgiXw9wMC9vcRTTRnYSLDgZTDEx2hR8d7nIyzMjH91n6zY
SGvo47qTZOxdjTVuDZ3RiM0boloKC6/ohMViOofHnvDb0o2NmyA8rfmeI+Wc4VGJ5+cUlqY4pkUH
0DQq3jgMdvX2w6AbGcAvRycQbLqSVQTDxjbhCjWRJND+q2lmEFnZgpf/0LjzIhyDgtMxeiOhPlKR
t0B/D2PwkhzMulMw3xK9DB1nhDgNolTrdZ6eKbk4hV+UBrRrQLpIreKSsZ/5CWFE6LtlncTKAEET
GtC3hrr4TH+Z8eUVp8wRfZGjdWRku8pnKao9Oq5w/WAKZDonHjb2T57JOFFfu1ESAi4Wa7MczFgS
t82WXEUQlcIt9s+F7Ke65F6+TVVyqMFzqeN9fP47037gCABUQGzQ5kdGK76I1bFv4d4oOIYHh/Ba
71NOWFU98eZJB6HRQ6piq4Fh8Sm/JvnBJGGAIEh1w0SBM6jRwoHTM3Tf+J0eqZx1lN/WaM3L9iaj
Bu/1xqIbpFgDwIhJd+6kPS6aq9zzDJoasJh9P8QLa8U6uqzV1URYVTmYZ/gexv1qVAEZZuPWzCo8
DTH/EVOw22V+elgWwEbWsRsD6iso7YeBha662l5sem3mIbKxVFRplhqs8YYw2oQ4Zlfqpj9N8f9i
8Rl/iWxPpVoA+oBzRQ0dpQerpzfy6EsyUksNs7S2g6QhNOltgseKuHtoth85bGSw9YDgl98BTrdz
vyKl1uORrRdnOd/lokk3qzEJICF6HWgGVrKpJf/ZE9p/NymnTzG+X7UPAP+GMo+YsnpP9Z1Zh0+4
s5J1wOIViic/0GE1U7otSdHLoZGi4WEYVE+QTCkaG7JkIvTmSGprSFzuogZwiuAGUhCmH5fhjDcV
xl3WvRzM/ZQTzifVOgFPl2wsX5Y1VUY+tbYgEIHArwc11lDFXVFABZCMddLk4G0iYfO88MZQO0RK
923+KGwMVNC8aNLnBEYyCIoZemCFrjF7buJL+KaRJSiEIrQL8ap1qNk/j6b5ndQeG+6uKaBjjng0
auAS/enD/t3p8YC7gM1YCc9cnwz6qDYcINA/n8QS0FneF05ONaKt0IWIpxBif0m0lvn73FvHA4GJ
K0fVlsR9T547Aqu0lGc/7tMuTcjlhaTaeogRFb1eHGhDmYsV2D/zUGLWYViSmIysC6bjtLbZpij8
PgvcMmaLb5fZrGDHB/etAnir7ZIj2Oroj+huTKINuvtRpA7S7ZhkaUh0/kR8UXnQfRQvu6V+/hns
x0KpB2AxBSKy8r/vWMYR2kAsvlmNr5vpoY38146WXGq3OO7vBKSPEp8M252HG1B3uC5wP8OtZ7wK
IHLC+MCsgottr2LYVWpfqysN5qjMdMFeHWrKsGSvYuuIQ3SR7e8AznRexs0ZBAWiMRpmfvyz/1Fj
W78yrpyx79u2u9tL3ZE7GMfZpVOskxbM1vejR5Ny2Yl1lny0S1qW3HITrqJYagAJMH8SuIOvK8Zp
Gl0lHmw7F05ACK9wxBdI4RfF2u03mZynUgdi8IboXEnYKwqTe6p11uwvytOFnKQ9xyjJTHAAe7nM
Uz2vwXrhHoW+UehNs1Q4jegj7fcdfXcqo5Z++Jtz1NvpoYQhsNxfKoWa8KXYW8Gh4a5Ky+YVN6pP
/cH/9Qqpcb0iWaPHdCZqepU4RR46c3+0Uje4MBCsOGiDPQp3br0hk1D7HZmL1q9cgewRJzRavOCh
W12x9otl6yxMmSs3pdDzK7/10RnV75Qws4a633LAxFXIwmDkw9fyw/7ApqR46qwSQDFQAZY+r8Bo
Uv4tntctLKgOfmA/GU3GndMBLwC/kV1AkCniY8SO5ho5MaClLXHCqBdXGAOI5rfWKXbn3L5rMsKT
kG6CJ4czvMPOMiF2GOzRY8phOd+oVeHoeZlfiIWBK0HQj+tFfTjgqvL2+zksyqlH5vnPBZoy7KXg
nwnFy4luPnBdvFw9gT2eI2eVt7rob86cm2FyZ4551LZ1SsWmCbQMcl22fr/eYVfD3B0guDW3i8Xe
E1KNO+Vti3zptyUHl85dLgPcVpvG39QwME2Ggr3YtyTiTAbcHMKLxOJKf3syuALvLulgytdc2Jrk
EYCHAL2InSlUyj2o/xj1zWQqfCJCk2yG8QR899sdQH/O9ySRpl1IZa7hdey2ABd2neyR0YLUyBes
RJyIpYWLs1/SvzQiDrOChQOlHz2UsWctvH/GQY8iHT7emza3eeVI1HdN67yAqox5wYogzNfDrcR3
83Ddd4UEn7BAwqwis4YW/0H7J98ubhpXjnR3cExp9zr77modLxt3ZKQC4jeMWvxTEnBsw084IFRM
AML1pLcEQZ7iBYvD8IC/oucfOGWFMD0GSMsh67FMXrL0goGgOXWwuva3PCNiwbSXDXoZrGt6ICLv
JBmlt1tgQ3voxSHvCdCWzz2LdKdrRYLFAhtxVE2PxLPJNNkg2+Us9XdcTra6mvrkEOWIuc2+CpVI
ZN2Jrp1390ozvL3mcn+5l1Bhyj/H2iRukgpzgQay4mcoBW9LswQ6W6Rc72WRoJO7mJHg6F46/d2g
/f+1mng9rzE+x65joHpSomSW7s+Nl1cRodEDvTS7iW9+pWn4j94E7mui4GOyHOSWTpgE0h1zpwhT
QVRi2wLzvqHFiyPSYPxQ22shy1rwtFn7lE17vCKcZLzCrip9RTpopZZOTDkRxIJEkLqH7mXtsqa0
mOqGeTRi6C2JMAMr5ldGhZAWEV8QepeXpdnWqJspjgXwhGidz01UhFIyMKAKUCRTAMIi67CeTYzG
nXD8GxdGwJNBB9d90SQIACfLCjhaa5+LiH1S7cxD7/t7PrifFgjsJV1kA55MGGFPzEwoK8ZNionV
gAij48wzvrSdXCAH5q9d7oICK5WcHGCFUdJU1SdMH+AdCNzqdgNhyLHd1rozDUUZzB9q1VXfvmPx
QI/SoalGLClzKUOCbPqixlI5CwUjNzDQ0XNBhHSYWV3Flor8/jXhI/JD1FTpNClaeO1v3nJAtGJ2
glwJATyCxIkvK4uBxmOZh7i0NOiJDZLqss+tj2Z4SZu6Jm+zwazBkSkQjkbAAeyyNOYPHbGsiJ4U
446zQHF6pjj4tW1cIIZKoIpAXK2qJDCVaqoaWFyG4lhsKTlF5kjVPqdvoUGQfeYQ4LUDRMqRZOAF
B9CdKxyVNDrJpb0TiP/qHWlwnnbaTMjNrnI+NF4Pl1Zr6VYOi5mG8op59H2Zh4cUEfkUXEgICn09
LjRysvzMXa2vzJRnIa/hN3gALBYHQmsq+jq24p/UNFmLAgN4v9OskHtqD2g47x1rLa8O3EpaHl4o
DI21ACNcpdTSy2Q0jBh2cd6+MGJgbPr5T2xyUaev7eqMRqLakLfZYGC4CiV/O5XrO+ct2kG2vK6C
rHQfBNONLwGsjUl3RREpJuLOcLpGoPLFdl/WbsSLLxCI5MRRMGfj4JHDRgNVhbnZhs/493QqgCso
SjRFYMn49vfkC9bMEJLGZz8Nmz8e7hxfBef6EY5xOEvS7axWSF4DSui6fFUR7vmlb7ge1R+paNng
FaWn6Qimp/Olyd7ELmvLhRj+oDupsdDfGPHZRFEtyYS4AuUUuW3UO7+NjZ5EVUxyiTrndH8rXPwM
mnZsQuU5IfK5+OoigeNra50S5Rm1H4czrokJqdEpgaUAcI5WsamFdKQtfPic89K5d6LDz5KJWEii
0L7MbdmpSUlJLTd0zZ3tKsp4qKre9wyekCtL994Jls/ZLS5+XUZTGoavoub8FW8wBjzYUiuvJXtk
td9KjXCiZPcHuqztfZlvDK1Hj1DFz8Vf26dxw9bbcOp+MJQAXpPcgILiHYUtWf9BS+jNMZsH03Yy
h28FFFzivx/jQmeH9hLtnoPgLXU6IKeU6RZQc4hHxdXBxMXt3ebjXsNc0dPh3wI6wtkpsh0WAgxh
DGUWL25fn7GC6dhvOnbEnh9k9wMzakdu+PiFNLzDFjvU8vOQlGTyzLwl8XzrUZG72pZU16yHDt2D
bMUKakDBE2hduUKXb/T5quk0DAT4/KKwD/Vlg3mbEzHGfu9NDzXyLLiw6eXSUJtPgHW7XpdnqV5C
mhVj1Y68+w9iCTo2rkmJcQPEH4IYZXDLWZ49S8Hi+k6l1c3WPy1K0OxyfajT1kyjB8yg2i1ZNDsE
7x8aFORepz95Sp23DqMOwABXCk3sjD2IWIsWRqNXcoZQrBCG+QQTEhq1x8W9QfFUJoMOLG/aoDrn
ZIwOBI//Nf+6R6B7+h+GAR+VvP7Vi75pPsdWYS3KXhEoAfoID8ggTzIaPxoec6FL8vyxBpgM+ATG
ft1RRBuI4hoHLQjKYV2XQX9wpnW/UF2N8KGbwqvCIfOOD4Rb2edPORJgs7b4M74sQhHYAS4JBMHd
lXlXtbfWnEiTCy4/yEvjiITGcgxeBgIEddSYKrbLQPbUWuwQaYH7+vYCeGTYlPaAME8mI8b8sm4W
tqMLhtFVjjlF3bj0E3Hmrb1tDNdDe01sYe/OOwq58H6POO8zRdEHBdpHL0wHhe+K92ozKomvMmWp
ewv3Vnp4fKkZaRmsiYJypkA5g+5dm+x/zMFXriDrM8FbCqvdX4xZrdfoaDQXTrO470WpUHrIwD8Z
fz1BtN+x6CAhoXeot/aKDXMDZO2EiD5bM+7g9EhBUZ3loi/VjSmyH98TpfCjDDFQKToUYxEPUIiY
WINSMRjUg5KlpIJWWc7eWnR3UqgbXUSxKwo72qs0gZTYgPmzD9xi6+OF+8px76bGMWUR6IAp7Okw
NEo4adK3cdP7b2n8Sm/lCqMZGC9SFh+0QcGFgiFvpc0NAOofz2121qE5CeJyVJVLW62Ec3REVo6A
dB1YTT/C+EsF++8rGJcLMZ4/Ums5VUX5wUtHhyi8cLGhDa6xx9RZ+U7lukIvhDeQKW76jYA1hx5F
GheLQX0HWhlkO66dcjNTxt3lXQvqwXrspSDHWcXgL4N88TvTXrYQSeLLw5vJ52qAxE4OlzZiqrgm
rGYHBONSED0ALD0WUhokrbc5XrAeRGHp8+LUcpjZ7JF2iz/6L7vQH1XQEApqkyjB4vXBSSeKnqc2
XIphubHtg7E22IorYrXyokFY+qViGTECZzeJZTwlUCqqU+9CUbZL1GRoydEymO4Cpuj0vCQjtGnt
TKkF7P6AESG5YzavMyGxk7JTLA7sAVpn9Vu4Yt2ikeGHIFtvZSDVd2+QUOSELDZ3UHPrFpYO3MDX
kBrfL+D3kmYt5Q/7NyIpwJU8+o+nQLmsbK63l51d3yuIfYGKHpqVUpCDy1P4i6BMH9EyZOwEkyCf
hiDMLmG9dCzs2dvqjuglbrhq4/Ffy6CE9MMUtkagnu2XTFHm1wTXYnb80Ig13heFXVxkfeTQ8jBb
017K4zAKlFIx5kTE8vC+UelN3bAvHc980MMGUKP4J9IA7neTomN3OCrOJ8c/iman1TmWkf77/r1k
wv0+aozjYAreNoyaDtXqLJbC6ADJjbxvuh2zJmrCZYfC5T8B7DrwYhFbAEjrvkA9FwcLBxw/akdO
MBUIa+1ugDHVJS+xa0kBPnosuslm/94w+vi9qxIEYmIIyeaoE5teM20+DobK38nX9z0JIC6UGqoz
R0eEOUaAdiE0kO2qToK2nfcv/42JKLVx912dIbnmuYr3bnelMB4gVhx3AW61kLbrJHFvi6SN069T
ZMIkBteexl2f9AcdPb1KgW1YQTfv11iVoCeHv4uxfbuGBFoU2+K5wtYX86nEOZ9iJ1iZ7qaoMWqy
hpcncav82fkXjq2whARMWv0hY/YUPkHrnA7dmqZjoBA6fYQ+JdfJow7CssTMhzdzKd9QhzAudcTO
1+1p9mYM2JGRY7fbEg5fdLfb6Rf6DuvUkfJMGQbj2djx+BQNjs8RwvL2IlNHckEdSzkKhqo1xBx3
EOKpzq0b2MeHc6sWbsNy1XY+U6dmqbPKsoJh1AmK9s7/IqMuMUjYPLNxSRWYyqfZqQHdJrbxxj9o
LKSR8iU3S3pMaX1VNRdlVNdQERryKl1wVXyt8oLBoyt+6XLtq/TuSjUOTJeN2Ca9nOzlIxjH5edu
O4rkfWKs4QxtQHi+sdmBkZGPgEau8Up24fFqrh7ry7SQJIm0fnYt77s42Fi0Mhm1dtWunfyZgK+S
HmI5qA1w5uVfZEPsl1kFDYL85/2xlIQqLwuAVTZLH3SP48avLsIHr2LdUu3aNyQWx/ZHOx67MppL
sb/DhWzVPHJMVlQexOz8oNR9SH6fYGd8gbonyqQGTtQg4KbV0OlqfXWcsKoMMpp3I2b9BnpAE8hy
TZM9jbCxf+s8ts5b5P82L7stzoTzjvbGi5kAiMtIq93sDD+5NYtiP0RaPiwAi1WRvyUStFoBtxyt
KU6LzZFojz4iV+dJ2y2x6PzIh80K8QnguCiCqH+Lc/QOUOOQ9976gZ3NJkUbzel1lEVReDr27fD8
sV5xyQtrJGSRt+zJFG4y8iTF2pNl5MAJeHkpyUPoWUmsOuDe5Gu2+Tj7wfLqoi6zVNX5xy14WbpH
xhlO4ed6JLz1gBmKwXJ09NZSQf3GvVZsox89FLFq+B/PyJv3Tu9NviwRA93RA7My71sez9J+dmDA
fAG4xb3ZhoKFiQJpbEYQfZm5UcCCyhNhlHFRap3xfLAm5ELW30Wnz79GvfxKoe4w5Yx1sVU6OpbY
ZSzGeX+UQJkry9QDRwRxZ2e00KbFb7/hCFA9BVUR2u7cjgnDKK8vUeaJA9P89Z/sfFCfVPcdh77B
A986/OpGtBFpuhMQ51WnVSbJpy+1q+iGzvUeH5fyt+8kYUhtvz6XnWGKuBdlM16xpRMb+YcIyEg2
NDszs8vCDhkeVZJ5w7QTqOsnFFPHBeQjDvPrgmg8q054HNDHCZZUbg6VQbV1Y2cWjUEYgOAGDgA/
pho0DRZBv9ZDbKFgI8eIH1lrBzqhG8iS/9C3d1IDEUiqLdb0EQOTW5lFzs+dpOqv933EHhQpCtoh
7wT+oq0RCR/sftaGwe5MbFYTw6WeQK5FcPudkpi9ojDW3kuElrCupVv2AHm3GjG+OC/v5enQHZMs
1bkLfzBRkPycNDjzaXTwKQhLtWtbAR/kfYymncud9JpevT8JeOQJtnYfA9Vzgu5Tk6NdY+28ZzGX
MGIq9LODq/S1TL5z/h6TfhaPGVb+kWHR3NrVTDoOEmRGi2VN8wfmLeO+Mkf2ecd02aXUKvdn3gOa
GfGrHeBgcU5j67pCWn1F3/S8uagma+L0YAZonAA5D2wYM3cyTk3W+yExwChQbIhP7wr5g9oyToZ2
9Rk84pEXPTDf23AkdhLr0IqOCN2RDXNz5+T9EQ5SAKcNp3TR+AKO4Z9NPqIIe8ur0RDRHoaVxNLo
hnC1sP+GI7BH58bY7gIH1eZAl9TLnmk87zfcqoZgzTp1R7wOaQknI1LFWN30sBoRcLFmd5pArNoT
OycgX2NnYo1rUrDpOvq3pFMo2Q7CL7OZlUxIdbx1P3tl2Xj5KbW+1wzWuyQYOVTPXV+Nww78hWBL
b5toZbIJEyIlIHiGKt3FLifOKY7o2t8eQJI6Rdnngh/rURCaM6JjF1rxQk0pwP3dVSvQLznYoifi
2xlB4ABTgGTNs+ENuzaOH6aSDTIYHCuaeYZHItttFpf1bPzVu9sn1VbejYVmzvhYL/MkEptI2972
oqRCzGgmJXpgcqwVaTRMmy3aXRJZq6JAfiVKJE3/qq05QLZ+rZZMvmprCWHnE/gzw3g00CkIhdwG
Azo1tTyIIZYo2Xj21svv4C3VgtA8diUn0xcwztaoIewMzIw+M6B6ChE7Lszq1qmkEF2jgAYHB4wf
SCOqyq6t8pvQPhtl1lIhwlTmRBkCWXPdV7bKT3+lDuDHeTD30m6B/GNe3m7M30h51573uPvK/Pkb
GYYF14kf78VHn/AdBpwBpHVs0inAFRKpY7dmFlgPLP79SmIw2JJBETeHK1wJpOH+p7v86B4LVXF9
9Wcr4KZN+U2nupkG4v2e3OonbWbF5LhbUELLyWJImYeKWm1s4nI9vyO9mRqg9SOjujPSHgeRDmCb
FM+/AXQ+zw3rqQ8ziFAdxfxDSHlXNPkqmLjImStCDjOGVe6Tky87mV54tJXahBCsxz462wk/3Xh7
DCLuUK3PJ+24jl7DxGi4zJLsjfvLCsgtCjGbYIpY1QQ4D+brjhBNzL8QGl7lG7H78U3iThK6C7Gw
GXZgooOZ9cmKHGONpvuQqdUcTeIl+nfXkWCfDnrB3RzHOcYkZW0gg9JfA12v4Uo8Or7qoKCMi+B9
zM51mqvn8jlo/w1budoWuHK/6CSiigSQOxMfG0JcobAil9RmfymPLwk/JkZiOrxs55aUiFow4b0K
H1EQyjJ26iSoIBDZNasxt6cSwg+ZRVb5MmGAxaxOfm4nq7JPkWUEgJYq4/Uwk7/CoaKk9fAJLTbn
YSBruEgo79FbTQE5xHJHv5zAjmHOPvgvq/ywtnJSEYi0EfyJLIRxtVvNaGyRwgc4i3hcTxT9IdPu
TtEHIfoq8KLo1+PzXpUL3T/sQfSF4Gc2DZE+atkslKN69HNuMWq2xMgc8X9U+VYhIoQGMhnX/P4Q
ovFCrnB2VAFnMKfZM0RyonM7BouRPCBWEWxsP+FMzlpcVOdRiVwztHLn+ZdFMsBJ4yBei547/noe
vYpT04VUSAwcoros+cGe8e2TwtT2remKFaZkEvpieLgfamVOr/0TAjAgiX7x0i0OOnhSk836vyeO
aKkZlViNkQUgyeQiqTuVxrk928MGBwAYkJpc83ZiGD9CAfrVb2jHBkoMhl3miX0SU6xNaqe90avL
Nz66qMAmuSuaU7GBMNEh5K+lSiSyORGuJwdSbx+VpRxjiQKN5z3uNBp/TIf6EGw/B5tmPQPWvcln
pSAVtUu4gASQOpuaTrBku994qyR4oyL9KPcp+tGazeUd1hshFHKxDOLzZNBn31hL9d/OmQ6ww1/O
za+ieT+4u30e1yb0VXUlf9e7bFhi5j9wqfBOarj7/C+fI5j5RA9Ry7PT6mDahdIxQyeoRCYSbA5E
jN/YVFAwEo+iPNSLJJwfDkWus3j0FBvSA94koUfFoC8RHe6N7Q5C26gsQIabGqYvsYUGonxBmS9h
L6MDGFCPDb8Tq/9/pvKmZrhtZ4UnDMrrl6Q/5eo96dlCOfNvYLWsPyXAcML+noqtlDNmcDXsNTKV
2/r8MpCjVMw2DO2QUDALfNZ3unqYapSZm8CuIAv+oVDlOPQWxJPBUGR0qFQdkHxZRogjenfphGpF
NTUQGzdOokSqJLWddjW7NgC0KCFOqyR9kMm93nXWNTmAhc19dmuzWhGm8xuxKrEFYR02+NTo+UdR
38ePZcp++SxcgAuWuLQ2uaxSygEtmj1a8CMk6Uwo3+BqlYGGu+qMrY/9tXvou7MUQxFa+pcvDLLM
hxr4+OM5Sswro8cKBf5LsZsw3pXzhhECaI3LHuBAMrkPBd87OhjKVURu6kieBcckdrgfzS+Sqljb
SjBvWijt7drvECLSiiRCxr4pCcOx4VRnn+wYVXpbjx2PqEjKlUiLdvuuEbp6Hcb42ODUUVWOYMtF
LC5NcI+UTJAwzKxhXVERnNwAy7VIJ02IubMgVV4kewfdSL14As+s8xsrI9WfnweogjYtq9AEhNkG
fU62GmCvH2KCwEx/E1L8nAyrdp0KrFTGLnh3oRHENhxPTx8enwHKLvrntkNbS3tX7ttPLxOXvnrH
IfOd3qgZ0hB70tqfRagzceirBNxBxFikqRdIt1onTbbsj2kpwivAqn27RK1PVcJO3+FgMtQeHhq/
4D5PiMUk5K1BiuJcAQHWSwrSJGCVjiX/BOXG64PSGMCJCsiA4YbYEtLnSbsH7u9h4o4qZU3Zo7L7
oC1w//5QDEyHyBXzJFaLew4RuuXr6+Pqf6CX9S18PZIw3u9TEyvApHUfphFrob38gQ6xt/uaXrQX
+QlTdRFklZJYYq+OuU7E7MGiFdmjg54mk7O363mUrtvUJZTlhW/WZWxpxXU/7JmG4LSVW7WjYU9S
HTCW6DFw4phqtznJHznqgkwTkWM0qk8E+TYQP2whujRSEt+J9cvrNSjqyQKqHpDR+pjmiozrKoUs
IfsB8AwUNmZcEgDsKkUISpkRqP4iZWmyHLU4n+x5rosLzh2h/wsZ1Di7repkUtMaZqEDHuAOuvqZ
16Wx0rGwupxISiLrxeK6i5CXFDOQOg+RTohugddGXTPG8H2sganJDRMv4ua6VKUBwdaZY19zBrMa
egSa5z47K6NKBwp3dqpjcRVZdZBosJksl+vfXE6bZ10r0gVH76n1WUj3lH5hZFF6OjxDfNkSrDeY
Vk69RN3B2oiAHbfYDrBsOSE1AqSe1BC5xIr6cWuLJDw224qymfrFuH1jQOiQE4gvUbT78bchYwNY
GZNWXSKw2uhQEPSJWEB4pjGmwUFaRp6CnRp3rm0K4eQgEXHMwhjHh4OmkSQABPwH4OtFLqjqYRqq
qlYuEn/HTCiKftMWkOWkA0xWzD+/ht3a+4kjmcPJmbiT22PxYHn4dlu1Za62PqCvbnAOHzQoOfiH
UAJ6wrZAlTEYLQBL91ggotbOIHX/3x1tEoKgLJMpJgB0rze7K4SPFGJa874su1wb9+0o6M6Eqo3P
97ZskJE/NWtjqNxTeD5CMvC4p2dXqH9nER5gphyIzsPalCqMDvWtJO4AUtfnuVAVExUOvlUuq3Tu
dMOqa6tB1BK9cRWvSOaTZ+wccOrRQ5qjaZ//wuypdctekHYGz0c3o1i4vqeafoTET5gb2ndh6S4x
9f6h9NWbMINFzaHCB9gm9oxeteL6mTy1VUVQEKggFEu2DzHX+4PsTqsRCmNaaReiYu3+MTR61Cns
oQ96G9wPJE37LcsSN/xmvkqSi3C6jartJNU4hHnXJ68UP+AmRGUHozxIP7GMHB87BjEjxjqAe0Dc
ZB/Xw4D8CoNGNNualdfRuO2UD+cfQP3XWK9KGb9kjDh8w8qPZEvWOYr5Jh1ocYuoDvgxuyeAH7RL
/CiE2lgKh9L7O7RUy9u7Ss5IkoP+nc96KTIoEbUk1Am2iPVhKJhQwiz7tgrC5sPyT/bQnn9KaGC8
W+NPEujabuP/+9kIzPFE6jrGrDTD5W7d0E8kcXSwxzBktd0+1rLvB/nmM4xmgSJUg5xZXcu9RIz4
8P5jUms7+hLHeE8SL7fqy6Oq0HVxuXbM5zNE6pnvI4u9VwdrzaxzBf+UNHjTYsmAfhhbB+fZsiKp
Hfa4MT9yIVD+tcKAXMuE8P+1yIx6pUTShZ+PRTaKfd+DQSqDXJQ5xgFNx7+WP1Inu2YprVHH0Bk/
87947N3DYtLjzNqvh+/YOL7sY7xqD3k4HOSi4QITAKB+HgTUpi8NE2pp3byWSJV466V1qhCgjq3I
tmaK1D7s5u4NatvrWo7RmoTpWeop0u9EMRde/Embs5GuA57dFb8MiW48Tn8leA75tmPUp4ujX63B
TM9C9vU+jGrFVV3Cpd0p1ybMdSVyXYnYHeodrNSR6Wjc034TmsgIgVtD7GwkVzN27LTPjOds4Bb1
w4ovSbcofLV1405Kf/upJXCA84/vsPbm4BV5Gf27nL9HKSVIRzJ1mK4JK9OZS2eI/aLbLxkpZF6Y
04Gd3i58B9dqGw/JSfjGeQ2L4ms/C3WDrJn3URBo86ELmU4LOZ/HmLEsOVhHOTiVSMK1ScWKS4jq
Qq9CL+6x/hQyfzZPf3otdRtd7ALOnSHNdOBfnZ7frzGM8uGT/mtkVlhM6rofCJIyu2ijPLYH+Z6H
w3hmWMCl18OPr6CTP8HEad23KJJi1hEm+2SIZ9DXVJvCr5vYxBSddl4Gk8lHU84ACE6gSFztn3XY
0TVOVXGis6/9O1BSCkqa6aWoS+n3sl9Md7osBxRJRP31KBvidRAAEvULLM0LIPeiQjoO8wNqIwZn
arCVDxvxgMN9hAI0Ck42tpE0kO9aU8c9I6rlgPl1gFaGHZt4urPbDzmVFgu1rD79lgRg03DAhBjP
+zuUS3Dr5XLM5+mnNvx7ojtuFHOmOAQDhUJiJqzziP6zP9yUs/PJao3+5/7AiCCrm1YOp2E/cZox
gYb7OJ3XXfdqj1JpzZYSC+p3ZpSGiMAaXRz1Ax1uG1lKRixzDHQutDPRiWPpXVMlRDPWx3NXK7qs
X4spwkwkEp73H6O56EKHYMEjMLtqWUThwJM0zkBvucgDhuQePYzgPp3mGrgFRnR4nBvQe9tTKyiY
cW10H9Uex8sBJ8J36e40zO3dCIvZRM9DfJpBhRZnEQUvLw4TVkL/WxxCdglHu1Th/ZXZ5z9TC4rI
RFpx1t79QiFKVqwFxjbMin1MVrkcS0ka1c8ykBD/pieZQpWTgllNi0T3EClniutjr6kTVhCYXY9V
fsmXzi7z91LXGX648JcQT6Uw2VzvyqxERddnOMDJgzEEuAxL+xFAlFAwieAYVlq27HNyQjAMmOnJ
S3/K9hpb/oAatuVDk8kMPoeYIcef+Dde/nu49dh7+ZV2VkxPfICoxK7lrLjMLyjBIGTmBJ46MiyN
KXm43Tjkpr3HfFnPPZqqhPiZFpRlZsGNDz5xuME3PThVitZRGrpLbNzM5cG6YRCclBOb1AoXa5It
/8BBYpyfEDGEU1mzGxA+VN2wQNXq5XuYBccfh4ritilleYzc7X1cLLzXLw2OYeHE8+KLr9rr0wC1
8KHFQ6nX7jCujP+Tx3y1A4gJbOJaE/vGFrBZkfKDPBgVl1VUCnGnMbBzOezWq3SOIc2+rZ8jWuqT
4CBCWfP7eLkq0NWSxS/6Jo/3xySkyOuocPWPDqbMQLrg2mqp6q1L9Jr2CzvxOwIESRN/ot+ssUaW
z1Pw2MtM4puJSlh5QTef3k+tmfbAlMECpC5lyJEdzyNhxO+rxKstkh1H/ABygCFz5sKe+oF/T1bt
B8S0P9cMoi1GgLRUMBrd1MmlfyyWNyo4qA+le8JNDHZ4TN1VJ3SekrdC+fY6lraOtWXmEo5UWdhX
NkifAtZ1Jq/ErHC8dXEsL4GbzgdOdjVePyKKSaANP60O7/hpKaEXfkyZrC1PoO7yd07tpnC10HKA
i+/lv8fK/A67w60HDz2oeyijvnGuSJO765T633vZCXQQyImmBcVBeBNwc748Qsr5Ib7P6S/mqS8F
DPLuEkkdzfs1Th6JaSsoaS62a2GsBH61O0zQeT6k3MyhVg/YEFocQLZ3no4MB8+RlcQcdacEjpR+
FqAUWZaqv95XwCUh328ZriDPxA86j6UJzfPGg8nWpw5fB8zdrIITDrGO/KPScgoF4oKNpoi+sXic
25YfSYEDFGSy7bX0Tp/7qCHg8CcXlj2UtMvQhwnIBJub8F1lV74u8H5KyiZ6UCUG08SlrpUTItN4
PsrQfMUjBCc6Ci4Z+0yCyHzoniamdFXelqD/9tzLfRr8usFn8WM57cWnYKZ6NAIguSYwvJyo8Y2P
A8xdCykLTWzRFMgLFyKT309mlHQ4gNYPKVCTiGQwKw82hUgxEm+ID0fLcA9yP299IqgBF4xp26qX
wGylENoDXQw3/GvfF7fuTeQZivDZFNEh7I5ebAoND+vQW4VNE8tHej7VcsRdolG9lvM8c+BoFO0M
Y1hSE0aa8YD409QqyijwK+ACHe9+QwHvaqlYXBbV+J8kdGN9pH4bz4YbbXDTwtYJw0xzZjHv3mpg
9dC7yJyH/QGKFFsf0pipqr7G8JrnpV3lo4o1bXqv49jg7Y3ewF9BGDV421cNbRy4uza8JSxRw0NB
l2H/CLdveK3iIqxrHc3E5CYzmoOEo/Sawck0ECLEGPBUxz2lSlboLasdTgrZqB3leVApF3Jy+LmP
/0rAeVo+dfpxaOfXZBu6XJ9Rmq7lOqRKQTUrrdaWqVejgWMTumRuhqKPvn1fUC76ZJShsU9E+gnC
ap3a++yEBRcYVSCiV7x2jX9LzF5xITC7T6GyBdm61csFxowDybSlGm84suhY9Bo2qn4pnOApd1Ji
LBNM8uBGH4lPf29HPwQIZN00SOqE6pNoS65nTtaHaFs3eXOWsI5mhlzG+6aGrUDM8nTgffCvZqiJ
slI1euE9S8yHG3ZIDuyZF1OcVu7p8NcOZHE9fKytumYMZGh0TCoEmCJisN9+6FTdsp/47teiFOaF
vV0zumhTU17E5I6T8VLNmTDQV4S//4i4GFIefZryvIJJCQZKxEB7rKwSnsIF44Oc3dMtdorF46VW
XWQTGcdNlZ+DGELXr1sY87e76pDJAYxSM0MXnyXPpo2d4+tXkAui7kuw/ZTbqZN+hjb68V0XEDoc
Uq3MDPWvT5s2qVy+y0JYOyZvDw0SBcA90XtD3/Y+5GORUdax/2ccHlLhCVO2JHN6tt3u4ACmIR6e
I3ER+pjgv96ktU/rFarAu70zklLHedHUnKTd9yVa5hogZ1fJXbRM8dQppYvekBHTHfsY8VTtgzrg
tcsyTfal3wmRBWIeT/0iZnBGYdCaVhJ2pp5S6UXLM594pRVl2byW9uhK74TadLGujIMycaSBXyRk
dhZX1W0oRihGbaFWkGLbE8+XA9qE0J6oi05UQ+4hSqbvhm90CxFNX+l6eBywnfx9jN22KUcnBIAT
zmFxh3jynQWZ7JM/Dd3kCUkY1c6J2KQBrVGjSjimVVwXruHYohO9svOXKFbLAzLZPrnxKGJgF+Vz
mtbtWzEgI1tH2tYKikIDK86SXr3RLpaAp85z9YSz2dVk/YTGIXPBc5x3l4JtUC16sLMi5Nuv7HzI
6Nvfm7QPcuTGAvPrwJ3HDgisXv8N66Ia5NKlhOGRoGaBMA8PtWmsElpdLlrmYhjNIwUjYn2gY0/k
QFkfE75mB6TWmZqbbu1aSyb9sto+YM5EcgrZh3MnS5zrQLzrOP4rEOVBY8nTCcyNBa/uU9HpVcsq
/DnwFZUUYizAwqJ9VaRNyvNC2fGOt3a6W0MGuQ/kZomeKntgT5mosWRK5LT5Vf0YJE0DOxarVP9w
P/FYyydNIqOBxwcu2pQSNdGUHgCFiCKvLKjZBeF9505nKs+uHbLb4NFEsw4mC8aZH0Ql8mbnxTyB
e8Vljj1bRaTwtqS4ab2cDOC4UqFYQzc2x9OAzCQNjPSk1DO+NHS62BpIR4/k35Mv5qXJDn7MFBuc
QZ2kkQeAip6HWOuFrJhV9gjybovJxCk4tOLNfGXKui5WacwwUngLSHuqC9QDmOiIXX9YuDxnPqKt
Rg21m+MaLMzQjh7HDj68Zz/y3JXJ61tluvkMringUxntO2ti6GTf2NrK0iTNlLcXNV2Coh4HWbeg
0agMR+OmH4Nmc73ivcfF3XjrRQimySW55yQeb0/MTpMV7FqSQTMP23/Sr5zNekzekVG9bejLJ4di
MbrIwM8XeMhWZWt+4ZC/vZDzTyvTjiCMfwqRiJM9TEFkchPlKmhFAh2tJLbczPBk3nwbNveCmrza
Wqq4LvX4fAh+c2Lw+7WtN8CEQUKZHTqFp5uC86kdArFPCc4mTUNqlOmEN5wekQa/xS5GDYpe5tfG
8sl74j9AOkJt+0paTvpq9+18C8B74iHLn6I/7lGjk/OH418JcqKaO40dZjgfyW4g7YpUF5/YK2un
1p1LDTRBld7KfwHdJgF6RzcV1J1ZT2cj+oAtuaXCkI2Pw1J7jb2NJ+D53hUhFNfJ28uYS0yxGtC4
pV9w1T995iSNYSugE/+wHdQuslwnxQnW+JuBWHJHcsOG0goNqF+TtzksvIl7O3epBlGCmMHlVhOh
lMy+w7YuLg54jcqCJnl43VgKaUXVc5odmu+98iUeQrufD/lemekAG+GmhRuxjUlWrUagTTHbaksZ
sFJiX9mJJu4fe50MRW5jU2SQq+U/hKVKNx+x2zJ6tMhyDIkZDAsEATu5Bu4kmrh+S3iXCPJ2Yvha
I5H/kThyyCCtrpnYMddw4rt969WVY/2l1nHYIpFgOzpBVOoS+wGcb7rEqBmeJw9XeuJEuAJ+IguX
LMNLaMLyrOyAx3ZokCJu5+g/56yxViMCqJBedlcX5lXKbqxaEYlASjA6Bm7EPLRYXy/FagrohtJb
rIQbCLJTsrZsSVUTZZa6PyA80wf7WGwwxMFHhG3atFQoRsiF87xtVVTjRb0ACNvlzFIkNGkEeUXA
jvfn1eK9vCnsi2VQhZW4GkRsCP2YvhJ3qeojgfs+m3ctC2n+uQnM6hM7MyDJGUzvEjY/YEy02dd4
YsZF1A6FwFwjKNSBU6iJU4aW8UgHLkw+AtoVxLHsF5aprM/q/eSxDLgnWBQa8uU66xuH81G89Xua
7Rvy2QpzoigzlUDpqBWU6ZJul5kgTxDIEGWZ33dXjhF6iDtrskJauuRwK5Dk8LKtxNzDqeSF2jWN
WbjRw5y9IbOBmVxCM3s60v1Z74DFVLOzhrF9CdsQOkrh+GUZljZxr69nCRLGpMuTfH2AzN2bMKx9
K0EIoD4pblilxsPjm/nAOSfzi/3tCn0YFpAOb3b2gt+4VIq3tFJqAh03caZcPyHzAFEbNoApVPxg
etIIVjFn9OHTtpDzJB3KegxtZqxl7T7vf/x6EAkP4D1oss+LKTrKKF2Oi7+ldevPTnnO5k6wF403
GjDTNqZtgmTm2tBkgWSNQ/iQTFupTvYgQ9peff/sZnAXpmpdtVluqL7cCmwlWtjDzCheRymMlEI8
0FEYHyZILLLhlqziYWGpG9AgHvnSw4SdP/PufwcqzpmOXDpjIRAODBuokQpsSF7B+/ShZXUGkXmR
3OUkqWoyi0VtP8+li4uBOpSGM19Lls7VBgYwm4BaQBCQZE3nCNBmwUEvVFIn96X7Rm8DIpVM/cru
zbj30a1JmF495Fi2IvJxkkk2f5R77q4i+LmLO6aOl8qjZlmuXMByT6JgkIa6XMxUXxC79GTWjNnP
d9oKak79OJfUlysoDDmHS4SrDCX+xRnIg9HVFJcout3L4I4zuhM+tuUcmzb8wUoyOqx6B9wLzpz3
F/KWVVEueytWN7cWu+3jPFCdiIG3L7f3AzfqQvCUYN7St3qOTIDIVCz5cZzhLgsEcPwt8qiz5E7J
AOBLi+cw0wb+T9Sc3kHh9bOL1fwxxNVrS7cPowK42DbISmyH4/KOJZF5qKh9ZKshrpP0wjzJB6x0
9p+tFXLBh/6nOw3vKtRRnAp2F1C5cGCClwaPcm6/8/cDVTMznbe1WguKJk20Ko8tsRza64dz4S7Y
iQI7abFXyngSSZxlZ4kuyWG+ealh8vR2Amz/M/xukQuaIaZZHPtjjXWtheLbvGe78TCyfCxYhdpY
ipOsV/xXgJcotjl1Ms4HIqZTbvGvYiy4qaYoDvKSBhRYVUiF666Be3DHDf5K5nSFYVq8mcob8fyV
ROnmqcdw93LSOARkbdsdj3lQF2LzbvrzfhzuHtI9T/It9HS+p6TYeKTwepCyASc3PffslrL7rDZe
Z+rffPJhOKohr2C8Y+bOIwwXoEmfLVQ6KRJJcZkanGxkGYNQVbrjoaMCs8KtRUWrD//VfcsI4qjv
QTOHBeGjV+9O3VzS2RYx5VZfnq57XJ98ORXNS5ETAa4Yn/roXqfK+RgKad3q0i01NThLCy47w/Is
bVh0NUayCK6EQVCndDdmqnOxpOUWx4SLGq3JQY7HGkSPYW0Eg6xuM1KjE81mxgv6OmCdwVEFsOrt
6O/76OpiOi+D3En9LUBrUmbGru3iJ3vEt0qRC2n6aEaJTay5vGp9zR/BBicX12Cj3klZxVu3uMtd
8iZBrFbdAteHZ/a8xsz8oUHNp7mD9XArLEQNfw2hNgqbjr8t0Rmsb0L+PdZZ+XkInS3f+HWwnMpj
rIJjVmWlKPfV63zPYwA8p8FHxXO4pfTMcvO6KFg429PFKLMSVdU4Q8azt8pOztoIHwFji7/hPf6Y
hptVbEs7FeNefuA6gC8gdb2DoP1IvyuAChQZHwxfbVwNkzT6ZoUlEPDIR6Bf9X9Q5/3fOzKEskpg
akNFxUmuN3Hr+E8aN1Z+DIVWRK3yjoWnTUaL57iZQG96g0FGlL7Dki+QTmAeq3wJm+XuDy9J+EHt
8DYN3S1qxf+IUjDV+RKa11jhtdZFqUGv0wDiZUzfAbsZR9mdoNh4cYtT8imE5TVq7ejfaAcins0a
jLKlEiIjO1tJHMDn2YGPbFyoMvdvGtzjT/MQOcDsXtqBQtuu+qVePn0WnvqVEpUvl3hN/JHaazJI
GO+kBPM3YBfIKT9YzSudm6i5oXD0Zjn8KTaPs0+i0l9+dVYg1ZBpD6sfCqW3Hsyph3jrLP9EsEHC
cFGZG9DRgoPhZJDE+jCdUJrCY7toD5o6sfsikQtcADhuZRSTj8ixyOLked9qKvKbJvIFvmCN2b21
tp8tKbrC9E4lTR1W6Tq/dBKtLzVHeaYZVCtDtE4KTdyFfC+ZhKWLFKEpusdtx3WSlKCFbEBdY3Ef
22GBdKU0LnOxmsifgTGsvcQQ9h9oXwdPZNOARX7oVOAVYccjC+0CQgyQyIrjt/UEh2LoV6RKOP7j
hzovFmjJ5u8l1eqE1aBYvzAjlgqRShTKh6pMmf4zO+bIDnEuF/SS2/jzEYbGFMI3mIcPtaonltkc
mkZhUDvkTLuIsY96ZnL6h3UxaeUrTCweV34/Rg9lgnhyHKMQI6gbZLcGeLV9wwlNrfkI34iycZP0
lwW+isTZA4VilylHHSEkq2kCJ06Qhw6w1e/HZg5wL7tudbjEhgh8MWY1FtF5cAEBzmJv4zoHZeMf
gsL83jHmtinhHlTX0pP5++ibaGbw6US2dECFIx8BUh+Y/AV9iZOCKoa0ZcvWFJAdFB6fv7K+kP8a
bYGrR4SO2G7ynhA1LmqgMR+a1/Ndm4gj5QrZ5lmCXHFOShk4uhX0DV8MPVNWfVAwj5nxzz/7jOV3
Ho/2uzdN7DrTXW/Iwc7c6I7WsaSnnNJ3Oh+wAQE/skZZIJYl+usrBiAHGnOF5N0wuIY88Z/MGv1z
EvJpoAZzossu3azAx0Rn4bdMGcyu3swzjD+eIht9vuotE5ATLk3SoRq1JdeZJ37ySkV3/HuWcQ6f
ax+WjEYagQFJ6yR0iuyP4plwlpqwk5/5OwVFTAZquI+KXxxoXUG4fsTJtCIcqHpK3D7J1Pkog5m7
wh5H/G5xxsRdNIfBVcpyKAGghs4yuHUd7z9b7o15BjHo101UejNNN2l3Vj4x0RnA8kd7QZszQjrY
eJMs/nydNdmK6KI/ECwAf7uCCs7NHScFsoGIcbd+3pnVpuvHCuK9zFnENvNC6wHhhTyQDjFjztmn
iiMCgEnyhXFw0D5MwvUI9JZCKNY2wwiGViaXiJEGMsRuOGnjwcx0JNpM8GuCZ05Bt9q5fdqOM5YG
QNLv3UKQM+vjXzcr+RqNGoGbbpwtqWeTJNCwOHeBWj3aWHHcqt6rERZj3qX+9+esbPL5gGxbmjwB
IbVVqOmA7Pa2mM9bu4XJs4o0mUfnn1yeES2fdarXpMn0bTyBy/HR2ny29r2UGM7AQxhxMLjIMBbV
M3wsn/ZnFDIQzxPfB7RhW/6IdDGzFe9hZVy6f1L2WpA83HAz3Irjdp9KSu1Zy5+paduUEXNWK8oq
6CkVPsuVl6XxitCrkeFKxu7e8XoWqCBmiU201DHKbrBEmHDQJTOWVJK0IT59/AIsleB/KQDhL0vs
1xVdu8SeeTx8dLBnwdOrvs2SXM5O47t7CvfAGYNMhPxRUs3saVbpdtPR6eQn/lKAc/W74fBs90Tv
t7bKokhX5dzMoZm6YzuB2qA2rLEp70yV2vp+/uHV0bJzCZxmnAnL/aSQG1gdcfNiTlLGjP3G1H+8
yzk2MkzYVg0V903xLxt8NLUngpMCvuaioaLFbtCsrM4yF6hoD22unamt0VbEjuG8Bisj2/pJY9I5
HwB0xbqIYMPeiqqqTBRhETIqlj3VeAy49tqgEkMiMMBLigI96UYdVxko/tyGkworuFy64kr5JGdb
gqJbkll5UMSilNU5QmmMLudH0eO9GmEqYp6IP4hgKgB+eP9V+ZYkGHaoCYYlJS7jNIre2EZ2Qz6M
bp6oolgrpmXTvhaypw6ObHh71ZkyUyxR/4zE8ycaBu3VbeHqnb0cXswaxiRCoeuS6KkcakbFKKz8
Xm7HVYsTUBJ7cQHgk2Dv2ZXLou+ioH2b1UpDgRj9z+vmtyNLwDkUhpr+TqiabMIR7tTGyIBLsH7u
AvQV1loFO5EqRIdAEwbb6yni7SOhQ8zQZZWRhT4LTPZ1XnD31JXdr6UGk7bYbvbful/3eD68i2x8
CMYVOivoeNoNa/2Gz4KDvdLXLlUvrQABQc9PIzaEAykwSF7xAQX6N577JKGECxQ6pjrcqpfugXob
1qxCWAPcbi+FuslH7Y+QdanmMJNo0bkfdlSvMK55BSU54uY9Z0pCcHUTgCGp71GyZSKYUyagCNDy
1Wvc4RBjWPyXYSzfWDLZCKMhUniGNLxOqQuG1rr4uGPIx2YiCpNX2H5E8S9sxOAKSyB4XvMesa2K
M168f0tv7vBQ8WRQ7mnWrHhBCRLrK3OlExINk7Ik1tGG1x6h+ykcWH1I/+mCoyJtirHTGoiXOq9J
Gzz4yHaWEKozyuwqiVyvNaY4Rfd3k6mAiW4VzqUkEx7U0P9tjXl6qfNM0+q9BbaezAb/41/hjFhD
DmgVINs3uvcRv7sVfglHB+nHbdW2db0NVPpQ7m4nFbLlMYwGL/adihRml4oiOnnRafc8V50IWu5S
JByY3ubG59vJwofPicRz4iJpjzL1Nx/DH4yX2NMD/qu2E0Uu4GqgFzMKz/Q/UthpFgnpKykPJzP9
xANAfMc7vSp8PQBWByGoxXTyLp4wWJLc4NlQzJK3TgpjnZ4uqjOfJ/sEWO4d/vU5fi+dLfz05PxB
qL3nitWrvkVFweknvP+SIqO5FOQKJTEKgsoNjDWJ6tKGUpArBFyW/5DQTjKehxT9KXXSPt+FWfMR
5tC8HniJ8KFTaZB3YrgLvOyOBT1ucfw73qR7Q/whtOMH3TyD/7zrUDlJUXLs5YnKnS8RhvPkKX68
9DfTvYCpkciwknsgc9fBwFqQSWPMPgnNgdTdKWzIUPaQqDLzLtSQ7MT/er7w8aiLYGXU3BQOZgF1
JIXmZEevE5KbO12J5JPMwi+CinMkGQY0uPMNSOZbKiwtdgMbeVk2W5GgL2VLpm+O7qhXXFzu4isx
pXez8XRfxis0C1uycQiE6f6x6E5NxhG98n4NKgrg7HQHrI3iu4oX8+i3sze+SmjYGBg/L/U/4BaC
XSGWswgTlKVDAOFPQQAt/Ri9zG09CnEgl1+CtqGk33t2qekMa0HelrGYWs6qcQ/6JA1JHGLS7S71
h61BfvCexWCTPB0JoYhxrIgdYcVSYs3PwyegZYEEXoqI5wio1c7gvDKIGX6cPOAz5LOm/OXbL8Hm
DjvmhufUHPEXmC6vkmGOrGbkaCmZqV7oxtrw9YlSq59JFb4QErhv0Z+cKDdbuf6Di4o0kdclsU74
LP/fyO1iehnLFd+QNDcTPgsjO8IgPR6pKSQYNsE6FWC1ZOV5NU1py1GI8FDoR8A81WsoEvWrTMNE
kNeSsIDJQ0pwTiP64PpV1neYT2iO6HVStne8p0Uked0WzVsSBdNJz8/sYzMsrMDRYo7HKHR0MBv1
06Mx36jzl4q4XkEtZa/6CbeVwllMuLHepilREAfl6lRd4F2RFxr2rh+KfPkRQgYxTlDKskiJmPMk
cOGCEPJkknmM+CyVASNi+Ef+GhRz042rsv85ZA//Qm1xHFdc5zyLHko1Onz3ur96JHPBSFfkFp/4
AOtCpSiZMsUrUFaEjpJ2WFF1s3bzXpfsYPEdB6CUttj2WI2r3ArnqGpUkSKqrqVzFi3nnYB7H+uw
1cwlxl2YgBWHq7yBTg88/9K2mvwhKaHGGt9QFlT/Jt+a93TNFK4IwE5wNRXN4Vp8oK5VzdX5OiMf
Xg8skOTX10PBOnC7VjW5vKIxTVbMDse5Cm1onPKjGmTZbeTcD1CLhiAxCGZwwIDNaJeUx/2/2E8q
i1LIVufmXJGTd1Hkx9vIoak4txO8lpSzq+gQ+HU+uKP4uQvSe5/Rc0Nk3Cc+ZWJi8cWFNzJbtpwO
hLUiOdMWWvVbqQFEmB9BiwCFaMrKoufYGlZ5CHRMU7cf0lC7eCjdgrWGHai+ApxwU9DJxb5eKMTO
tNUIblALNSKSDgxWnT+OlLlG81k8VBHFkLu00cHUeawKjqvDgpdouZWez0dsvEomx6T6LecFauD9
R+XYF4MVU7zyI3AsfmRm7i2pFZkdzNmOl8Dhq9LRL49IsWv+zcCtbVEpr1RieH/brkqQJcWzyK6+
PzapMY3BrGA97sSfgj6Oo3kXN5y4lxgcMSjz6aK7ryCTD/YnkW+Rt/btNCp7Crms9I+Oxct8ViC6
WhKJUtV2xaIeYPHgJ35eeu2lWcu/AZnfyBcniSHql+ilLJwojElCVgz1ALeIwARnhRgBC1Q18H+l
szMvVIToHIKP+njGc1FvPXJf51QOOL8+dPQ9IOY0230xJ8406adHHUevL+g/qERnK40XJKz/o8QI
1DoXof5b2/Ld9ezDE5N/FaRQVbo1lbR0wcJoIG/GxRDce9no+T7nrt0UlhlnDkl/Uq/qCuzBAwS0
OXycjM8Sde270B1vYKadjQg9VyaubiJQqfJGV8mgl4nyKVpAK+trsFay3r6J6sOn/sa5hgpgw2Qh
z11DEWgZBhn0vNXARXn1iPmkZ2svAA45tpq1gjrIoZ5Y2WmRzT/VjdVXzD9RVAE11Sq/e2VUa/cn
exgC0CaQwctqoin5QbujK8KUl/NA3j0XMmGCUEvmvx/6GPZwRr4hSTNPRvH5m4XJ4B9c5oQ/EZzv
KRjBIsE6qLm0mQaEVMFZNb3YpU7imGakwnLSkFB3Qe+2MpV6KG5Vhi9RFyAfsaVAfBmQ+SR+2rQN
szSu+ZjhwvHxt4NbQxn3WmueA/vKMRwu27fvRB1L5J7OgajtHji8LdIDvOfOsCMadY3NxqpnKhHI
ttHLbT58O3VLa456tDld3dJx32/jTd59Wc24j6Ix2ohj2hzXlvHs+e8frKBElK7YKRqKcqoNvrsh
hzWXACI+k/gU160s5FSdFuxVEWwluDaSsCat/1nO74xrUkGNfgRioUra8UBVQk1BasqHD3XTNPws
b8EitNxwcCH/O4RGrVcSrtQk6g1WvoYurVQtUuyqlH9e5MktA68k4JmM8L6TcftH5adJ54Ddasxc
bBTXlpcaq8osQSMq/eTDrHVN9h8W/xa5X3GRZlLIGFU7uqEKZaolNXGWthb6WY6srCbNWJKwKEtV
/PFheXws8th0sdgADm025tOT9vPuo6V+CDu6xyHkTkAJBFP+xTcQMTRV9SAbVocez+TycCYeeuxf
jQ3MITdBwYt91bxtcHh8qF2+IDaIokHPcJrnqAxqmsykZezWrkAZkUVtFJzNM1JNzsG4VKIm4oJq
z0/x34GULeDBG46b2nJT5WIPcbtf3HnONIO+6s9tq4yUTFONGKUoVFXMGJrubdjsKNlaQksh0ka2
TJo0VnjbPZhFN7ucNLkd9rbubaTwJ38Tp5lfAqdslbIsp7zMYZX3WvPzOlzqF3K5PZ9AiRYqL48M
epyreiOfZt6VNFDFn5zm2fs+rJJXYI/+Fox+rTScsTo51OHOgw23j3hQ9SOp2q8K7f0Q2XZ6yDDR
qpn6fP1Xeb5jrfXNYxNDWNVMcmu2kLD8NNpkaZlRkyz4GcFQcLf3H0oZPia83a8Jj3TNX1bXH766
5er4H8P4UiRS6/wq6rW7XFwAMA09wKUi+OM0eKu1Ik7yfiOmqDRuv/sBuBK8bmaMGHt6yeuAnGDi
3Zv/Lzhrka4HokeTdP9P46q8MZQ8jSlTowhQcN11+dSqfGBANodOSPPOzWbotycMif5WyG5uIMXX
ZT3cCn6xC+BUqgipBQtYpRpl6rWfU+r6YreSYOKZxWVRMih4PII2f2+0+rvN4SsTvtTvss3Nxftb
sQGyR/a90IwBeLovMYXLvM6T1jwKPMM26Mj7XolKEE0rv5sr3BtBmNEjI/aurtLqObqlzHBwmRLa
JIvLiK2QLX7PvCNNr0c2hmP9zuzSz5AWi9Tg4fRiVNioqWT7JIJAwQOQfoDltPsGEedShcrA5S2B
9MQ83N06m4+fRRwQplCacM/oceKg1YcAEZg1FaYWQpV1xl2bYvUwpL6CKR3z5o2aRA4YqTI3KPzU
1JKe/bOcpz0NZxFlYmJY0PHK9Yyo0nDaPsZIqp0T4F7tm+M48FFXUqBRNxkwcMNVsPZ6hbwZqft0
LEIgz6PIvTRLYFy85ppOBtZAXAghddvWnA==
`protect end_protected
