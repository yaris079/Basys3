`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
W9OZ33fX1mh62EfjLHpW2JpPal2vKe+HyjChULbWsn6SCOXxspCzTIl81L5u7Yhl2LLY0zd1w9Ss
lCFNf5QdFg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nWkKh4PxKnlizRMnSVczSG+s7omR5nHpNq4He11trZCi0N5WH6F30cOimGjZNhvPmfgIfnGeV7A5
4jBOwnW8C6nBDxk/NJS4T+vQpaaPvCjct2UnF/KPKIVr/GEPCFGjyC2pUxg3BVe4IX17c5Sefh2R
KDaEFCJ6A1XJd5v//lE=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V1sO+xbQU6lp1HrNn+zh8pXZnGbPmd0TqWCRVKg9Ir75hLgJv7sejL6QtqeaJKwnbe4qjfT66fig
o6D7EMs3aW+jy6WHaHvUdp1ZM3S/X5EZVSctQnrAlnpS2kujiEU3OmJGqMh0aAlxcRELgjzrCyWQ
0bfjdzabt5k+q0SHxsKzVGZ10aHKSgz/YY2DsC3JErX8gw4f4TV4p2902ldcCGp9MYaAAem7dXcK
DdB0rUpcCMWfvxQE37rp3gNdpZNFIJLx/uwZCpZKZKz7sZzf7ZbVYLa5D8/zO2+ohvPBqsnqRwCP
Uh7k2JHKoig4kxA4mRPnsLyXh04BbRDkwnuZPw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
z8v2qCZDHpydUX0cdWLZ8ywlx1Q7BcGgUbPq/1MDtQqs56+eaLQKH4uwIHEvfcvm9LxbTFJvhc/T
c7UBM3ILv1QUO1dQqGc4QJ+eiWpdkEXhJrrCVwSVDbYrjvYCWZohx+WjLYY3JkikgfwgYhkPhnJq
9UtPb0CMA8PUoEUNZbU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sjExqRm8K8ILfg+3pzRc5ctb0k7CHJRbWgToIgxkt0el5xOzdj+Ku8xoCdoHTrxqAAzdZ67Ivpxa
N607XrwiZVFRZ25xTUgT6pGVCBGpc1HOZnbsUeUMxj/U5zu1iBuqIFmPazAknOagG38xvOpUA24L
4hYNMcdkS7ttu5nykP2h1Osv9vuHRJC7a6O4MdJ2Sjbn+fFN9QQcNtNnnm2WDfuVGX3XVKU2NQAa
+ZTvERr+KzF7Tqai+o7zmy0Kr+DxPvXikp+INaDsqThLlVv1fEqu3LihJM20Juumm7qg0tdwjnuK
CHQbdAlVVFe11Chdge2hgJMTusCjOtZ33uB3Lw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11152)
`protect data_block
yiX7X5ws70kqOjp6jERU0J4KtbH+YdXSkbZnYYJq8v8gtvesLbgJuRV1qnv6TwZ+yZmfrFIIGva7
TsqCQduPEch5NbuCWRtUMqVQKTO05TQqwhW+ofjPgDmJH4BV/GFP2002qfZsTOeWFfHaKts5Zyd5
cr/9k6lXxyktMu78ft3LfRvSMXV1wQ5pxkcfRy0XdPIiut1368PwP3M9AtvzM3irEij7SrunyBay
6JIc9ZA3j6ep2lyrXq851mvLAa0TCGh24jKgWxVMzfYy9Eo4K20bIURTnWzN9bAo/jDmuakmvYaQ
vJzuVeqaybg33aw5wI3mY/nUqFkChypVRVBNQ71MMSNvKkeRliGrO6jvD8hjUNONGdJQ/H741iRy
MHdpj+BbuoAuVhNq4/VgVSC491RiYEOT1SXU4He2sFqHyEoiCkUCU7y8DcgJMNa6fN+2fSlndBIf
wHmvukwyGuLskREuAhIw6gSaRCu1njHuR4HblS+G5g/KXmulXmKG2YkIVmfquzPtZFkCrE+wpnzH
OS82ef5O4Vi7SkQPwiIkR/jklDqpukHMyQjnietJSWwLClBe92V2/BT5YsFNVoC6Etz9emreFI68
aW12sGwLuH7Au4fUrZE/b+I3JQLtn/EBvoWTgMotphm5OGaadPH9EoRNdO7RYDJnMbjgD6pAgy2h
+s9/h0mUIKeWZvrbxwR0sxWVFMmc19KEqPyokh6EIGQOVO/X+T5toDj/BxVFZqSpUTkw5R/6cIZy
orfnc7+B2gmI1Ut4a8BUaWo8nKWT9Yqx96Rx8cW9C89hljnAwkdCOt5tnkO3gP5QG5Uo8PEqLTCN
um94Dby3BzZFGZelDUwbpdoXRJ02Dw0ThJIlHEyrENkcjwfbG/LkIuwUuvajEQdMY+bEzhiKQ9ku
cCKnSgqfTbbDANk/R87xnRR70TlPhajV3c/T9bzdp8w9gAWYNSOxeztxl+HOB5Wm85QC4VWSkSHQ
5wpt/CU1hvJa+XH4j1Hs/fn3v1Z3BSGDOf+RBAaOZoAxVqvRZ2hxEMOpEWoqqzgd/xCJ1MDa0S+U
rjQxJqpVcubTl05tcQMzyyWjxqOXv8c+Urmn9uj7x5yB3r1WE6aI4K9YlZeI1iJuZOxqgbUlt7xG
DinklmLBHPoklGAl5o/H/yYlOU+PjxUpf6N8FDxhUlGG0fCOSRKnqxAuvPzlSpGopKIdg0fU0Pli
Xll+NaMZGwwXQ3OAzWa4FvT9+FQe61/chOtsBO6KVMggFVgdn2XEQ9lVOdShd9FAIIYfeE/k8BTX
bTeGm8Zm6bX7BFep75rqzqJ/pHPkw8N7Q4JrtW8263783jLfgD2KHkPBEBs3WfL46i9KL3ogLMqJ
VbljA4infG83gDdInRdfYSfitXnhL6EGfrJQ30QvoqoGmFJfYTuwsV+F9iOcf3V2uTLME22YhsD1
GtYi88Gc+1L+FzCmHpBa+1zH1t/rQDHcLOSKhUz3sZEWxV3ILr4lJBJ2HkKkq5KJBpjhACafL4Wf
5+UyqKTikAcgGt2WbRKwVPfzPttT/p5KWZACiEc84v3R6vTEh8rx1bSrXiL6JXvMvQ8x7u+kDLxL
5CWmn9LxNUtkPdY+2eY1k5RrHPgpL77boJwgwbb2XRbGxKI6XPoJnJ9nHQsL3Lw+7KFh+ydjZoon
RTtDe89C4xucaCpALMyBhQXYE6hRT3EaJhBxudRnWviNtk+3UoJe5/DaVf1ysICtNNB4hVXhWSQZ
sDSxeemdXKJ1sS90LqdjP/uWXiZlLQEFcThFCf9LOch6gegwStbY6s2frg+EUN1I6hBNaitzdYD6
Xq5nUVNDOTZGraH2wv0HQaE3R8DutCoSh842OOmMEw2MjPQNFZuwzoQzWfVGAlkF0Rn43YMY4p2h
ZQAdKSoUjEfDBY+Fqphx0edT6MHebg1CICNoSdl1HhWtOkKjrph9fUETH7lbJEk6HxGtG6OiiLBE
1HpEtD1e0NIKGwlobIak/lCCPUWjkXX3oLaX8TxLbWvmP99IC6sYlt3QTHO2SeIexzLY5Zzt+fHZ
Zdt9YuDrnbb/0/OnFn1E+Sx6RqqLNE1xX/X6Jfjg8LGX8bJaFrkB55j2b2EVksPKHr4mwTvVKpFo
4tKWzghdgxHcfdLBylRM2e6tXta8fl9WAaTZg8Ne8rkfxsc4gmppByFMzWGVdHnuRNBZhgB3jo29
ceQ3FARFbeQp7FS56teyoryePDhuxmpARDdB7FPCveNcg6+pp56pZap1hREYyIbvBIjbER0s4Ram
1+o8g+nlMMCtZPl1sfBihXwdc7paFIIKECChxKqDD9v6paAYrs5ZrZjTlHNI7fSXkzZd+MzBkGnV
aogumWZu1lI1w3bJKvkuzEC0vFeFcBdywUNJfRki2LSojS+cw7jFztyM1md28RRqozyDAxQRoDlG
gOf+qzt45NhTdrs7wJaCsFDgZ30rJDMdTk0kbN7vrWfDXjBmDg0pQJw+4fhBz1bfWk31E/D3Z3U+
O71yIz5pPFNfQ6Dw6AYKTeBNCmkby2zfubGuMbeMExlu385WsgiEs7ReiY6+jXwSufhkMyebn9Ii
vvN0m2B3cC4WLbU7aLhTVFXfePL8xMMrNguR3S5EAW9Yi9yCXDQMDfdLe2/zXEPFlyFAQKPgl6zs
mYMzYAIuNGzn0yElpa5T4ejomHod5T1RcKrzOj4RvAo+ZZgVkDdPFRVT+lJLOT8hHOeKkSKUmcWg
hQH0+6gbNAEwaH4A1YoEZpOLMwtebn/irzoLqMeJEqfu1ZZ/lMp6mz6ZO14vemkMujaUNOPjaP1h
98g/Lt9rzW6zp/fzS5EHL4FauMh8fRVInkiR9Qhv2wJplVQ9vFGM3M55DVT0VX02z9Shb06YghVt
Scsh+4VP3wIwLFJFnUb/NGSx4cLq1wI/VkQj+UGJYxDjhvAgijepPmcZFYC84qj5Zj/cn+0M37cy
asSU860BYKxw3k1gq1XQz7toP0bIS8maAXAiySgJPQfxL8xKyDA3Gs0wnjBqQCWPFs4kQYqXEXyj
2quwzKw+cPMcb/eJfg2A9/8uMYKQoWYHAeeFosU3I03zPAVkrqlcJbdWCm1YyUzTqEkjteVo4A2y
JiXMKR/NqapuHurLk1hJjrZNXE3Vw8NMVacLkyfqYp5D9H9zecQRaQ0fL9EtFxkDV856Q/kz9Uyb
2N0bsFPgNyhe/feNFwcn0PAunbSncC8InxLwMoxGsTfRe6S/T+wV7DHCHa6R4vSnrSVcaY4woW9M
hEs2Z7NHHDJCJJ9i5PtnEBLekfUCQiuXCodKnx1hmcXbXR73ZLhtVBKMWLRZmt+X+Zm41bgHVotD
46a37PnA8y3oxHFCtEWUo4UZicjAEqwZGwlHbHFAJVvX2p3CcJdPDwYZMJdemdNeR+wscRZXTg5Z
plmkTD1ghAXTLHGMhG0eqlNdbkJBjG4+9vISf5Y0eUwiM1A3aHq/01GO62C+7WR1vHeeA3cbwB4W
HY4F45YB+OilY44e2XNnckCrRDVO829/PGBodHYGVgEXuHFFXv9yp0j42BhekLzA/BYVyZ6J8Kmc
WMon30axEwchwU/7cpMCycqfgB4SFOV0VXGCwqCLvXNebgoKgXp4z84OeEf8mqZByRXZKGt5Nm4N
Qkkj8CnVfWCho94pfnS5Eb3oHA23izbvWLOKBOR2Ulmf5m6TnjAEnQNohC6nlb48tQ7/NoTQBozY
vUaoyyIk2+yNBpx9HDdweQX2Jy8vaiXtETGZYHgf/nSPw4QT0hopOCSXgLXZHWAa/s500NoWQJDj
HUTHrDKt7WowWCs8j5Nli4E50Bzitk4/0qz2O6l2fmD9SryLGLjEKqdRRNrndEFaRX9m9yR4bwZs
p4YZva6iNQzU9Yt0v1JSbvKpmPvjN4jz75EmJg9VKumc+B4wEopKRZ44hr9M5olaAw8bJgOcfsOs
2l7wC52tgyqynTSSyaj/O67IMwtKDyi/9S5mGl4nxIUiH6/fpJldDXIDvIGYjiqKuTvC978M60WN
ZmKXe9sbR5yH03EkZWmjVNBV8GJAZFZew010cRfwIdvG06cwkFrAJb/wxjTCdwxUtmCjklycb/1f
uhkhc8xQtkHSoZuvIfvVu1WqMNpZckae6uB99a+Vwfz1qNoAMrN0YZKvzylGtRZfftaRRnXRGgYV
WmlEt4L8XtwsJYeEHLLr82Ngzhh886iXeAyOnec5G0oMmlLN65N+LNuCHs9dShwiUA53ABupIzfS
pPGCoG+l2FE4Kw3D06lxVJDHoN6IEJP9J/bt//VbR2IAtrj87+jwJrGz0jodrFTeRHYWkGrcEXrD
fQN1rqKIE1gCmDI83zYbVLX0lv7Cw1RFnm+xktiG/dHmfXUEnP2AKfFsZMcbHIn1vkN1UwjCVyWx
Qy2lM2lPlqjMPGc5q1a0CNS4H99UZtwNn5zP4dkbB47ehScO/42L4gS4nA6EI2ognIyLBcnmrqE+
nQFsodGAO5Ad2UuNiyFoD2bRIycAipICRl71Znd0zf4YR7k6YObKadIuXgmVWOb2klRCkTmzPhA+
1X17QZ3q8VLomdzbil86wMopG9zN4q6oDDLRayZzJfCYQMbByJW0k2U6KcJVv57OlUPo0vd9dRyW
OYDIKq/9kTxDEuu5igLmlC9nWIR8SHPeaTDdbarOhdzJ4C1d7BcydQxYuqT13QoR9OIhBz8gahYc
5MQ/hJlTv4yP3eMeh0XhcrB/eOUKJYIRu4/RgRL5skynvNyLxf45FW3ac18U57q3Zr36Wep9hqPp
WPIYxJ6lbiSg29l8UhXMhTOiY3YnOLVEBeXA3iHJ1h5oyveljF44NHQIxYZxMermudhpVp0/dL3C
sWDbTepbdlrDlNMEkzLS9Ztn4RgsXTVTYjPR8qqwhyMwtwb0ZSRiWafZ6xLwC3AycE1IBYcuH/fc
C9fCA8fOnVarHjj/DMa4VRaneY8tcmbSYUdXr/Rj2MAyFe9U48mPH4R6mEHqBjyQgrm9ZRwOAUSE
R3JAYsp4JhWSSG1hcZo2K/Mj7HtT1Lgxyo7RhkGIX2F5YJz9/c+tmhSLm/hHT7XarBbaPcjmqzPT
xCR2yyFpWbHdwy/IpAfu3o/2cGjJoisulu/PewJ1yBRazclVIZjj9e89e/kRYeyUNoqY556jCOEr
rdXI/Q7bsqy67CobfbcWiNxIpRQ5EzqAJpPd+5dHXWXgu0Vw/gHIolD8DuTqkqlW9MPNbTVFksR5
wV6n5ZdDzO4IxTRjY6pEIf/osY9wOgERfCKW4AhbBxIJNbN4tr28cVU9Yedp22lgIVNBFiSzML3j
YggmNilR5pU1a4XJ/eGh6i16VmNL2zrOhT0B0dRjgFTpvCxTRy09CuQsr7lCE6XmvY+yrPzZJzBT
rZAOstfqOgSqJ7epETY8ly3fo9IQ+Nv3UoDr3YnxHz6o3Ymts7LyXw4QrsjuMi3JBOf75NQnlPtH
jc5oftxPBKWxWR2qiN1kUTkdmFik8bjGUPGDDvNRAWuK/FIl74Nynw/jwXpArMFvJZiIzUyTPtVO
oJqqgIEvc4L0pCxyRchG7IX9aIOCqZ3ShvoGhki015wmpX08UB5tZKfkfX9InA/HtM5sdpEzURK7
9l5TWgwj4yOTBNr4un4Ap90sz9CMYUb6DNEfq5yAHyiZMjpYPV2YQNBukWKRfI8v3Kfu0zHbVZD5
uRiO3M9ennXIP3r0Qe1YvLAPz+Dt0yzSzcxf4ZweGrzaod+a6TM58P/JBWixoK1Kq7nF90UtLlfe
LaZig0bNP8jRplDadoy+MeZ32KyijtloRDQAxm/uh6gYcXw/pQc3SI7ZSPXbxPLoV1ZC0tU52fcx
MlEsn6qSPJojU7A9XaHqW2V9LugOCId9+BJ9WDF5y/SzZbXs+cszH77EGqcaaEFJO1Y7Ma/SOQbS
ohctrlUtJroLAL+Ol9I+HfPa21LvDxHTIBcAMLtI5MT5GhobPyX5P2fBD+USxEjZVHKnwr3BzpKu
LeRwOhzPkQ5ZZae123cz9ExQm5m4uaFs4icM0A2hqrAht14H7dbxgJa0R85wDTZw08R2wStesdV2
W2of8xWT6j97mvwP99blRv/z3jsivkzdNyRwOh/nrTZS2G8Um7b+9/iWR5rYA+EJT7WJ8s5mCDGx
sEaICUk/755eu1zPvoL8LiUd9LejtA6+BchDlAL944L5tAe1hC8OCNlKIG3C3vFMc3jxn3ewcoYy
uFP+yuQNprUTIFOLf+/GpF6ychgTX4JEO+D63jhe8Fr6ENjLLKmDVLZbDejGcfkvFi31WiXGfJ13
PCwLtuceMxlYqxPEpuXj6pX3r+OX4RA1Ex/LjxE3v8lP+g703+GQUqWuggn/QdzjzmovO74h95gZ
yVk2KB0hFa2/vqI9AXHhq7aA1mTtadIqCKVd7K+7tAv4UhsNDVrQpBKD52hOEsTEjbq01bjFGR32
cr+yclHcE/1QKJnQiEsilId+emxQJRGpPPdpa0fjJ6HXhcW1YKGRka0ottxozY0jgEnaVrGxjdTK
2U+iB4Nz9DTkpAAB0qD4QIDOhvmiXhOzRTmnnpw7L113GTTuicryUmaXoeQdXzh5oXfAIJMe+OU6
wwLYVpyDYSkVIlwd+N+O+ioLoqqWmSJ22ZgrQOAJmk6slseStYjzziTkPF2raTtKa0n77upxBwol
GMoNsWrF+YbaQ5q17+qnjCDTIkZMtdsRUlFO5mYddKfcLVgnDK8jlptfg37Hp0CT6hGhmuInkxNU
JPFRYoIndH9bvJtrcsrHDWkyzoDpSqrR41GpLcbEqyAsto+dVBo/NiDTXrdha3pWv3qutJa0r39T
3rVNXIntLzulvwG7JQZMFPry8CeX5igQUJSfND6+TZUok0S/HeMRuAW0Mdd46u31hpgPBKoYIZ3e
UeVw/qHhsiHl52dr0wyqNAJS8FmMZNVD7GUedu3DYM9hAeD/VPsIo+08dWHGjvy/dCSMTgO6hvUZ
mGCcVTga8j7VvLo9gNvk3PxAQLVsBOLOsOPnWq+gB771/+3DRP5cfMDFCfEv4N3JCBug8XECrQyP
lG4O84P5Jbmyd7tHlofn9M7ACMabbcVsrtUjbYWQZ/LCIIUHXwjjSYvk5T38Dk62DCM3dYHf4Dco
0rB1XRq3U0YftNBOA0W1BpToVp0CvD9AoYpsFTq6Llu+sUVqF5ucsuyBtlVAL877TP+yzOWxy4iU
uQGC3VxIVh3RCe2I+PqnbHdqDDO/UJT3EbtqHRtjKME2ZZsmU7TFVScv2o5UXStDCNYOA+CgbHdi
zyTa6D538dYv7uCjERvHhIKmH8pxj+LIPX/7WXXOIy2t9Wz8HhrFH09iXkPoDiD+iHLLWn7ZMhv7
fWUZHU4hEDxuvGhvkS3+Yu39Lucy8CzO4mcX26Qzun4KTPdj2Fy/4mepxtz15HeFQZDqagzxNzSQ
2jgHhsYhhvtK3NAN6mu3HlYOnh4aB3hmruIBD5gOqZ2Jdi6q4HOLEXUSmIIlkddu24kEjZCgxOMF
1Myyl77mBc3p0ZWNBicN6AfEwjLl1B7MoikJODugXX8UhLem9sh56b58NFX9ztOnZWal/KYDyel+
C3KIX0xeEfe29nhtvMaIe/ZAZ+E80WiRGCtN3W8sgxXR3qa7wE3haqHXBJ1bRIcty+G0sKD9R6iI
dQycwo2cUP+/q12yaXBOTDYkmtRYfsp1nutR1BimHO1Jr5cQr+U/34r4P0Q02QvR+TZ4XoNOuCgt
dEDa2GpSSKz7y/eVBOoKIzDhG0m8dQSGawB5PKqaBbK/MZAd6w5ilVB/CSIzUZ+P2WAqX7GOdhDK
2iFzKDHbkxRKOtpygQGJxsVgyrLCH8BkC7Uhq6tSEg5FV1tcbbHD6ZwDwKp4wvH4mWzNXFVz84XX
UN5fLeoYfayp38QNW2NhS3JSzRJjaXcVOdx+OHx5gtwz+S1d3y5wOCNFSB4I94kWDpPVqr7CXp1C
QpKzC8xntE7KsaXXz3UCKtzlqhgA5qEnKkuW9qN7odHMLqjKncer9hAzLHPXPBygL+NeeQo+Xirk
Nx1GgryeaMV44S6rAjPFu7nHuy9x92xmA297377YueW5u/yhCkPcMFnyvAUOSp+tflo9tQffHLRD
s/j5qyZcGD1NplqOnZdnoTRHTenVr8f5ZZZBOGpK7PRtI/K9P+3eQRgkgC62cT3fJbKOnw1Cw26y
SJsUaQD+k2AjVOL8pNWQxLq3el+lw6eHvKaLsH7ZEiGEDx5ly5+qEdg88CF27nt0/uJaMqsZSkMm
Bj+mRHhW64asotvKAoOC5o8GF5jhvlwz/9vakYO9Nq2oHmFtrPu36vZum+jedvFupzu77ejTNBFb
uUXZH57085+ZNX6OdF+rEr3Y9fdyNo2+mEf/GqP9v/E3x+Fprlx0B08JMLbcOOj/U3jZGSeXuJcE
t8q2X8gwBpJF48/J0vlmwL3/sfI7I/XNwXKpa8xnZmitQVkGCk7HC0AwVFrcWsG8jGytqdvEyVNs
Mn/o3PbWp11fJfWTbC2duticXx7l6pV2R2zcepsldZqMOnzVoQjiDTJ/EusqWu3JmTWAzGayIE+F
hXgoP5KYspDDw5ki1kLziOq1WfusZZgGqa2xrYygqLl1hOz01HxZ+ePJfNRrY2HJIOP1oijdnshh
aeQMGhlK1bmE8osC0VOGfSjTymrEnNi8fqPbb4o9kz+2VbwNnmQSeAvu3itf8afhVQWAo37xPA9p
fqKK/LYQnUjGeYVtYbr12h22JpoZy2pk2APT4ooUdxFTv1BZ7ZZLLEMTdW8HdyE/auMwWTByzNbT
exkjQun5GXl48JgXUwjtfqnb0MhbW4tfuV+BZNije2C/+LOwcDiiChYvofkld0DyAKxcBxcv9Kmt
xVFA33+cfEZOiF8uYLKzuP5WjMdG/ZVugJMZ1XpaXPc7kcQN+CeHWB6vpkHm9x01Der2z/3iKnzk
Sq+sfyc2MyLw6Z2c4uNrEMDkZhw4lE2zobqVP1/PfALdgpCaDnnPmLlLRKW/8dGTrrmkZXt6WY+Q
8mxkptwpDrw69XAvA+vTbLWTOeVgNn76B3DBc/rBNuo47L1urCza0ydJmjVV5rSar4viO4KU9Pf0
kju/onOFkHysdQOoXxf/qpOzDjF/1zGF28vC2aP0VOQOuspyyrBcuz41fqnIhGs5VDtgeDyZ6jiI
PLqUgmE8NBoR4xFtDJx01uXwf5fFwiFaZo4DLoB3q87nH+MhpcSu70RygOH2jxykYY6lzmuuZSrR
3SmdLQ3F12Sqpf6ns0oC/vvmbT9oNW//HXjbYd1Dyt9PF7FWRpfFG3dtWog7zUaZTilxbiSTXGBN
GWFCSZWM8fR6myb5T37lNlSyK/d3DL95EvZwUD2UGZtRbQOuuUSQgwFMem34rvMXqv5ykx0zDuK1
yjTmyPqJ4zLMW5blzKZWzFyXPPQ13u3QFrnZmHnEm9hIETVXS8scvNRcFc7QOxHHN95uB1T4jNVW
qKxJUAC8E3Dma1QL3gw/g79XIoav8W7j8438TfMms7IqtuH1q65KhS3rjX7+LQbSXiTNnaXlVmCT
NvOYdEZ0TalxvutunIEXHbPJZKds/eppWg6cQRHByBhiVlOqKAqwLiPkd0NolnTgQjG0UZZNirHZ
Fz/H0d8lm64z19VX47hTolJV3Gcchf/Ru/n2wF//vnm7lluJUCDg+lQQyCig5utN2RGhE4Hdwkwx
NR/7SBNaor43VAAaCKkrwbh/+nPe/A6tb//8kmibVZ7MpfcJrSYeDDNxcPmdJOwpmfYkY6tKIJbs
tpNDF9cFZMvjDaQvyP8G8kwUi3Y2ft8xA+6DGqban8GTh+EpU0fMTUx5XLv3fT02QPPFBUvwjuvo
tuz3Mo5CDaEvu1dpdLd1klbvjN21ifoO/JbFfKnYY9kFHi8ISH0ukXOlReoBuS8B0+DZ2A9cfAr4
ZyoEU942zBKXgD7UZXQ5oAcmUMHN/+qrR9BiL8ZtLbTK2LWjqEadERiFWDm9yIXhGOqr7uQW5WJx
w2JsLWofWZKC8v+hRwZq/LF+vFJ+UC6c5qbUpRBv1PtXXQ3AKiIWI7Ed6YrsiX4ePsd41CIV5LGY
Tb2tM8ifEnc5gGlw0rHUi08BGVvmBCQOukCaNmF9KuUhCHOkRw67Czo8GDMEp/NPoycKfV6trSbZ
B7UXg5idYEwwWbLA/Gywwm1UYkvzehsyrLwQfMKL+hwX2P9zOkIKunXKEEDcKgVHDMCzEAwnWoIk
uTXkA8kU4aC3feUVNFGWQJkCHf4zytow+reHEmuDfdxRW3f6vWdASkiZeZh8qIqZJjwQAjAoz7VB
jhpBNG/QVJ6Hfd77dyF8B/MjKZjX1e9H0qqXQ2NEzxSvDfho2Un4IOHluKklU+e/CSKYihrvLfSj
I4QpWKRNsFdpkPndK3FCT4QjjCLEIHwmvXP4Mj9drbMOC0wVCT0hDgqVumolGf2PgAbAmvS5K1qZ
v1vdZRduHOzP9oQgQbrGiIWbtZKVQI0m9KeKmZmcZpdB0KsRGZte3HVOTWYLMhiH8RQLnjoZ3pxg
YosfixrBhrHxHuJ8Rwz42OGzsEfSUZblE1k7xQ3S29dnofGwozizixwBzwQRmxyNl2KQZMsmh3mU
WGbDtu0lHb4LmGR4/BveIWcD7okSBLo8P7fBwDsVJ1bvRkQcIkFIrc+XkBgbq0a2EVrDWMvkcQ0x
HaiTrwSKncwGv2r6nPDXqWcqZNPoTIEy3KOSeVHYQ6ZpIiLNLzhgm8nh6BabYRwwz5b3I9oCsz1V
1xpmDWuj9Gh3WUVxe644E3TaGF9PapQt8z5L6UVD5Y0mkfsy3qkwTBrydpvUWbEJA9aTy/rcRPvl
FSKA143So61/2lfW65lUTBNI1bLy67WPadXoGT8OYJ6nwSJqAafogTWUJ+204nawvp6o9WXOitR4
w9f23jbJkhLlBc5sB8KnMGvnS4QB5qwqGv99S7P/y40+9pK7Ql9WrZ7zffbn5BkSxnmfYIAiHwaB
jMbi7tifZByVmFW3d6GapxWEmXm5y/MKxASdoCLq/FN0EHRbFaKL+sfIlBC5M10tPCYmTFweSxQe
G771olYCyxSZnhMzuqmGvOGHfR7G69ZizWUU1RuUztQQIyEO9RIV0q2oNs/h2rkyDfdMlCNsS7QM
tklTToQRiJklu6Vxjfbcuu1yOasoStjsYpXNcVrsT+x/6MHQc/GXxTfN67z7hjn/vkPNfikNuq1E
V6PvoT+OgpuMbdXnd5DuKWLxdqyb75dC2MYQBNEiMOGVgB9x5xjzX+DqmY9rO6fjWwa0VE5+yItQ
6Mw0HA7JKMvU0mu+zzjdjMor/z62k5uMUrntvbVp4kKmNslvKIoViNUM6bQHo2UdOVcrlKhc3Eu+
ZepJLbi6mkPKxYqu9/TN9DWMxk3JHmWWEi4Gcmt1lXE0w87QXQZSkLJOBElUgfbu6pNuiOJ1TeQw
VrWjPemg4F5sjLtwz0os1QeX9MGTZP9yF5yuDdeqKNh1Zvfe3pqVg+svQq5Ltz+ZpDbqYSfGc4OS
5pzW+HNKO2YdKyXmBzeahNkjnibOY9+R6gQqUG20a2AZoqFmgZaKaoH3uznY81qwL/gORs6TcCuk
A/FTqEh7mvVoBdCXLqpEsOjZHPGmrmYnkuICA7+U8IcQpHJWAAMh46BylqvkGkvVExNKv+ZM5tGO
0OZ91AcGOxJfv9uQ9B8LkERPfeTCL8e4u7zwPvvYzUXziyNkMBja7zjzmLQqLVp0C8EFg+jASNmo
mwsnXrRbAAQvoBLaoyssyK44G7u6st7utsUxRhF3dUXLc997jLqvN6vyB5MhjbC25IKHlNUXOTHT
jqAyjy5ne/9qFQWDZKtyYxxJtnX89yJ96JOi2FFeMKXnl/1+ZVbT1PQbX3BWAyJvEjO/HQzWwXIa
JsmdqVlyKgrW2+977/KhflwofL7ozkBnOclbXq+p7QI6Xo59yd6bOoB41YqF76S418ZX4BFmNiqt
Dz3BPs8U4MfiCWO169yYx6cQHZpb2E/xdUkxrkjEYfLZNHG8QV8Mr3ZK4aNWEVMsrJKk+lYJiOhd
aEEHaMOniUy6vGqyjaYWJ67+uwYB8cbopeB6+yyfOj3oah21TDio16qGtNY0qPxvwPzukfB/hQBS
B8Px+33LWTDdGoAjeUw5gHMM/w++K4sYDSVTdgeoUhzLy84AF4rZ89b1Y37d1HcoK8nqUiP9pOAO
VJmK8WjXt3zcQLa4ZvFtVB2L4YK18ttpz8F/TFuCeRBMnHT95lCJxOaHnZ0RAL/VwFk1ApoHQREX
k294tKS3Zb2P5iqTC8+JqCa9bG6kT/hDct57+CI0erLV56jEnGA+UfT6KuA6MJt/Wv8thuWg6bsg
tQW2bp0rrll+SQTyqvy32pURIFvcKhqCISlm3GU2VsAZm4/zmWoxo1Ck/BwKFtt9q4N6gMQwpyzV
fzaY3hQNdnj5s6OQajCtbUdfb86o6EysOLTXgkj2wgbIbBruLybGMU7zp8ws2PoxFaqtP7PWJWrK
a+C3Lyspp88yPdvMYEUIbEMFLBEPqY37xxAswM+pj0RYLCg3n5++h9Iw/Bz89CF9FJmB/xDUiFpT
16VED5IVgicQKZvcyMEKawmjU8u9RXaL3uykTEAE2Bkfsu3rlYlfqbspY9MyVx+23vWvIxUL7aze
gmz/FlmwKt03pqFKZhjTPg4rS3Neb5cT1Bm/2/jKqhFter75TvIyDnnH8ro1V+OGJ1PNHRQJNG6X
o08CFhjXEm3/enhDN3lSvzPmYT0Zn58c9f0ZjwucZ2usM/q7A6dHzLBFMZx7FvagcjiKN3a11Z4d
D5ZYc4be1PbZK/s3xG66cGe8JnReJ2T0kcjtuTGfi4oh4BI+vmGPoUcbs5RGGTBB0OSpDfDortZh
Tlnuqj33If9qOPC4O1GumgwgPeeCRIvqcsXg8IWGwjLhA+ky0LTMCa8C1gfxm+vI5HMIS8fQ1511
IIXwfUq9znfAvcmvre2UawRE2KkZBqvC542afS8JNpAssRQX7++R7vKTI9QSSBc0A1MZ59zg7Iym
G63TFmog8Icf+xLI6ugQA/S4ofpiaHhCvRrdL8sntg+Dwe1RU4WRMeDaWK6SIapn3D982kDeZRGj
vJmRPqxCQ+Bz1QpdTBF1zX3IRz2AnhMMWxs8ip9BwQyOXCMs4MwUPOqG/j/cntUuGTLOPHVtoWmm
+MpML2AnBFH2gW3irG1QoN0JzbWlXL0rKA1T/1rWsVmToFsLiZr9iL/Bt8k/94Xlo7VDXWOCMQZN
vVmdv3Yy0HJwdYkPxp0DminfTdjtkwTuxTtbR6CiHnV6BMuTNHxDmb6Q6qzPZw8OJnTzIUmy9ag8
of66OGcMOXMczHp5aM8V97r96yCUmMv5DwS843r+dHJTGLgN3bHDuRbqLn3umcwAZdkurl8gt5j8
er5I3DfHjSgbs+4fZbKiYQyd+wEZ/DCvdXvj0XajDJjcnrU7FIwRhXd8J5g9mQcYgcDQy2IPJuDy
1rAnrY0vnZGu+TciA20QZAqmNCOIHoLQItCATLGPvVcoDs++HenkjjdS7lEea/YtMeza/6yh5uYL
8zxaNZ89cNKRZKTSIaHPVfgnkQwfx0cLLGYcbKTtGkQFwaT2zHiBZxrEh+DG66/rBp6PleQvzFx3
R3nsO5vd+zMQz9VzHI3XLVjSeAcq79ie4YPEAwxhsrw8uedetHKBoXvblo9DRV3PuCq1t8FD4ssF
hz6ro3Y2iEAjMWCIq8VvZGhD+X8nkWUEa6/Wp6DKTS7dsHLjzeoSsYeYRdSEp/M1tLiu2JIU4KPM
qMNG+JTNkYYArI8AAB5EsOGpuJzrQEARrke37r8kkf7lkdXel431i1Q3UZX/BuKjyedy4SBkKH8/
IisA0A7r0/VIgu59BEFA7s85ZDtJVyjNb7XG57C/5fFGv+GsKjSM3CSsjY5RCh3Opwjzwy+raGmy
OXsP4MKyAsiUUlVvUauxS5IpWrlr5DxDjdM25ao0mPOCyhJJKhD97dh9UQaFh4yqEVKGMvHz1t27
nwdoEzp2/+yiPKtXYyK/0y2pP1+FJN3uTRXdR7+l/YVv1VOqbpBB2WECglkUHf3oZ6lQZiAQI2NM
n2GesTBgmyfVqR6wo/fSFWpL3X48fT6Rq0fmXMRMGOe6Gd5LSj/yGVYStesnMFpXF1kd6Cz1gC/S
fP5lJBW95cUGAx9olX15gy6+DypqX0lg6Gu18bPPBiCSTjl3jraAAxuG7DD1FIf4aqGLV+ouCEpd
vj8kErJwmO/6VW0u7KvNLNy+31Tyopge5h+1YNRkJou/SjkacEiI67Aj8J+z7IO8KNloSgGpxnt2
EFQDDzEYcmsK+6Vo6km/M61yBCk1U2tNqWRdDtwgnWFn74bvQ5diC1sYjG8sbi4ZIHTpwnRsairJ
sjRNs+4Vqg+oHjHh3WqtIL7y/hI4H0OrfdwEkKWLOf2fKBzhidQgaC+cqctMlb0fLAAGvIB1AUkt
Mc59TBIJ2/FFR3GQ9cbc1OAUhcBy85wgffWLwe1DDjECxcPIl1Wbi2P1E0L0bJ/REHZiKzhWdaS3
fcnDzFZr0sk1r2FWivbuP3QsLu/sSoDQljl6BWgjtZvAxA+lPERUXonFfwG3PxHa/nkf9rHAw2h/
XFVffb70bC51Z5LXSWkwwkcGruA/7FBkf4Z8WWuY4BTIfjmEUNJomxTFh5JTnFHP24iobsXB0735
oIQ5nBkvLYf7Icdh3j43Vkwx1cEqESQg4JQhJe9NMwYtcKqlrv4r3/MEcRp7LYRLui0NrCjoAJQd
lGEQJaJcLY+f12HmEH+UUVzYc2/y06rNdeamHQzAVlqyf6G+OA==
`protect end_protected
