`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oM9evIXQkd7HcYtdMAyQ/pzMuJrixOOoMEkn7GeUeMug+eUWXAY0jMb98m8uNGVn+jdi5lHS5V5V
9nhzY1B0LQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QBzNK6GkbfR6REVaWKnLyIj2T+DLOzlOHcxNXVZyGh+CLDlqK/7/2/el5fDCUfMmWl99BS/ttOLA
7rdQdKZsVSYp87vpl7p+RoTnfBGTOYynyFWzHTEbxNnWDWiHwkSQ8PJjIpMFVzG8mJTUvXsTwfsn
haS9ZgZpEVy5+qAOLTU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rKD6QumD69GDkqEWnDkt1q/6wJSzYNZAfusXHRdunGLapBiz5VqDea0E+0xJMUTy00kBDMc0hdR1
kw7PHy7JMdtgvHW8K40D2T7OT5sKOK8m4jgt0k81NECeV3fWWOnAe+uePyHjCj6dxGLqOMa0XKro
Nd/NumAXyoNWqfWNAxF/3wWuOM6ZuQhXmCoItj+TpSsLGGROiN+qaXM0wg6gu2+16k91rXwtHjXU
f3JEKZlUSKp+Y4F9r/E1bTlfH36yJXclOmKj04m4hrU8INDB+ZHaCvrCgFzTokD9uTPbcvGcgeWY
CoYi5wd6nd1cLUjVEX4PVfKJye9oMdTa3HD7ww==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Vxya9P3UpMLKK+DGCitP57WoIjkpNik+yUA2J28y9OqEAdK26heW6PMnwmHBmuuemnf+9x1lJf3b
3Vn5nJ4afTAqby7Vq6huy5M+xaQOb7qSEnpFVkgyBl/Pu/X+B/wg5GtnUOtXjXXToQUODMnYkr3z
xiIAL9KCJRzHAWSMmDY=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MqovIAo5zvI5HNiUKMCVgEh4jEGdcYJjSeof/Ct36e1ilX0QHcIuWCa/ZimNMg3d0NDpSprUCU3j
WwoZqwBCuxTsv3UmLb96x0T3VJycyQkkcZWF+iMxPzOR8ptW3CjB6vgo9H3tTy9Zj2NmoPhLBfQq
J3/ZMo8oAhv54j1BEZtJEqwc1xnIF8ceEuwVasLJqvlvLWI+NNzmc/Ju9ZlTLQ9iBaE6qY75TOq8
napv0nntp1EGqfoge26U7ADKlLd3WTogZPdCWwZ78TtoV483HNQFhHjqbeLTqXQK0oBPGPWfYFop
PxwEKl4ftUSKTmv3LXf5vrUCAAnvnKWU7nRRBA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7328)
`protect data_block
c/2kKoUp+1hSznCIVocjdhnAH7lGTcKLpiTMuPHWngdwniv0xh8D2imKhdG9PstSZ+2a7Pw2L5Ui
Vp70/FuibSlFhzOT30tWPJXct3onPPTkLBHJ5lo4PDSvryiCeAm7VM8Tl5/HtJ9qqSNjkGRD/rpX
nmHCWMf5PvGd6QBjJoKnrj9fLsxyMlcFJVAZqLPyedE6jnfFVx9tcRIoU+xPOE4AlLcjdta4BM6U
qFYINp44kKk/OT1uP/0pycodz21z34coWEnZnyhhzgzl0GqAN5RwKJZ0fngspkc5bXv7jAZgSR0O
nLdMiFwzlwpC8IgTxEOBp5SIoXJp62MXo6FjMu6kJDFJHvd6I3XUMN1SK0+rYAUuX63UGAeaVkMJ
N0IK4gN/pHMnNAMcorIDS+IqNYhYtmz80HY5jOksKc+ljuU8Z7lAECOsAQdaj6psECcXt7wIdnQ0
p8LseRmeKllrDgYS6PEi9lvDA/0lXzuevBtfItnX04TyrToGZzD8vjcWmAmyclzJUsZvyVKiBzYU
MKuJ73Oh3QH+ylJzHfNs0noHBCZ0JeQRcWvcdSCQRs1A9n6P+M8MVGvRBkJif1Jp85rKpQi0IMdY
gxBdrezzXRNf0vgJ76buTrIKE5xownLvx1IH94TjaAwx2MOlOxlf98dA4s8hEgR/f6suG7oI+ank
NxcrGj559pvDigVeqhZ9roWTSiLGvOrOv/4wokMVJuLVHeXG5A4U0zCdD4aysJR4s4TUGaqSBQWg
UHTQQhdSX87ffg0mZQdJ8wRIblOShgBagw8/eEQ2rSmUxQH3BWPAQUhTHx3rjg1AIK4/uoRPIda9
3mhV+EnuPZP+db3tuGTV0+agC8KSvR/UPWENcXioqNgHKjxOTJpcPmyx4NAr9OULTZvUlDA5C8X4
rCodsK/pMQDsL6dHcAZuSSHHXzgDIr3KL2RLRIUqe0oRQV0XnDbW5gsaaOoXdKjF6ofFxwTdqVs/
sEO/tPDwUTpwj7MupeksiTXVBJJO1qaeuqZ3hEwA1+igHmXZKO8cDkanRTm+Em7zVAE5GucQnb5V
lT3pBiifeke6ukP0Nw7vjDEZ+geMxIE2eqPKrJU3SVMJnR2IDv/2n+V5IgSfQeBg+PHJNvffHX6p
2lDDzzdeaogWmgzH+CvsSsGL/fuY5JyOYtDk0JKd5F9fBfnu0+T37q6X70Eik6zzJn6bC884yQRr
3iO1KNgvi8h3oj1XQU01S3/8UfiT2mvreMq2UUrK1N256yKHZao/lqLHF253LpL0+Whf4/bYRh4H
Q/BzCZb7sjp2dYfXc3N3DGd0+c6aUdsfzHt5RbKqC7I2VfoP2tYzgH0lvkI2mTaj5G/MAqO2jmQL
5yM6LVJZY6mlPksRYds0iZW+R9Z8SF7YX4y76ho6lKs/Ai/ffs6AiBL8A2tOF58Z/ET95XgZilQd
sJEKpMgPH4o7YTuaqRC52+GeTlXjU4R5yq/smSOOq6Ih0Ua4fbTId3jvnkJ26HW4lHbVnkt5tA8D
2MMpuxSqW7h5xEqb/nUkGkgnMo1EWr3yx8MoL9M5/j1/J9EBZUKcQJWJeMrL2ZxKgiIhOA8TaVEc
paF+fz5SamJyf67zeOpR/ccKFi6S5l439GOaK6lKFiYU7vfoFyg4rmAYeQZf3JVz3IghpGiBfXIS
2coeMs6RgN3A4d0S/TKbeG1aJhGCm4GQEbG9TxAwKS9eylUeEPheYXA9i1gXsIL5iu64rS0+9mH7
IQ43RiQRkBgQmzDueyaZM5v+j5ilhFCVCYxK1rpcOID8hONBLOEYi/4snyziW2GwoQUK+xbS5e6/
WtqFvFNBt3EvGDEu/hJAzEVegRVRq0vWkz6pr06Osk6/bmZ1TLHp7iEduNHS28HWtDG3s0zNktRX
sM3PWKSBYnguNKL046uV9i3bRY1dbnyQjgdtI15CX/pi4sLoar5DB+IoG/Uv1DLh0n8yep5f7bJX
xsNJRbgtNhxLAxdgRvgGTS2Pd6ooznnrtvWgUH1TSYazdr++lg16YInG+ySrrgqGWTYM+dO6+tLR
fvfOdo42mRBesE+oV9E/yUeXkVydhfHP2LNoVmik1g9IRdZR/IhkzrEsFqU3PBBKkvd1z/6Ua91f
5o+3OU1zoyw+Z61XAwtrXX9xyFXLQvstp1c3CPk6SSJkBLi27zoVBLkYQxb4LqPtKTV3/j4WKE6g
cRLH8ouKE2a06d9m3c/vleex3q59vGl2yOnNadzTwFIfVkyosTrkykzIaH0cgW3WBPUW3nSv36FS
Q0Gn6tIPeW3+qYwYutPY6zPVeuFdUeusScCkU1SsV2OBfSI7I4RhjufDJ0lzMGlXDCi9dr/fn/bc
W+Jqjht5uJ+Q+Jl8N+RFCNeUJ+eWHUV5Gnm2r0TVDQj6x306T1aLjWiKwWAOqSJLShP8u5ka5oYR
A1Ak8cSqxfyjUW/aLYVDB4/FBozlC1lN+eUHUno2cz8yzTLEZl6JFewIs71sV0KxpoW1O8Ohsu/3
jweaun5k/+sfI8vWcGFKdGTzbcqZaTZhjXJzM6dnyGrNhUoQnt1GIUcnDeDY1vx69ML4Vzts/eZq
0qxCJ+FEjHGg7I/+C4YE28y6TaQ7SQv4JU3OGicsZXdOtg9NHFgD4u7LgnBYWoEKsS2BjcLRgr9i
WQWWVXmAFQX5sbiij9/bOHYkX2gCpO791fvd8tabVhSkqZK7+eU6TtkslYcr8tSVtA5dOZl2s/Xz
9UO8/QalnoIh+rFIprxbTtw8zSILCZesV3OrCDneI3dxHQ2a1JMx/8DNb23M0WR29r16/el2u/62
5NeRHG8CibLv1+gCKZwwo2KK1IiptufBOMbt+vA87s1X9C4uA2JrSQpS2/C27mI3F27ZDgR8n9zR
w0WNJdSFWnF7jEg7VGZAp7/E/2eT/u92MXZadvhzfxuGJbHmpaXq/Jq/B3c0SLIQOsY6hEvrq0xC
xHZ/Lj78i6GuNV1NABUnAhnKz/qL/T2/dUG+Y1kGq+q7CxmAysy1G1khJfMfZCdnIUXmX5EXRoRG
rAaqUHT/VC/lUDXWjharXKzSOFDPnfWMLlC/RNKeGzwr+Dz0vn4w1S3HhAKV/FsNZ1at+n2B5J79
yJqVvW9SOyXqG8zQf+GukByclkmjZ6rSMVPJ5T1dlsnq78SDmF9KzBSIGadBz5POOplwkG+/u0xR
FWH8nup7F7xux3VK2csO2TOyUyE3crxo3v4FQKGV7yZzKY+NDJDa1sRW1Hv2aMpK2QeQeywV2Y0R
k7R0TNcK/CEnd6qOFjRyr8oCatgHiGen40Rw80brjccAfLSZlM41APhFuyV07poB8jBkqEKk4q17
Ir+h7+FsGBaxTF4bpwJkN56nmrfHNyGeljUjYniLwpsQbGf3USxQ1HwO1xInX4mbdz3jkmqC7Ein
Qj66EqnYMr+wnWUU9Nh77SgaaMgHyFUTOelXSwmSVe1/zFYb3VTQwixQsR12oB0HDrKt/zNVF4rI
NT6JGnmtQ+v6fQWG9rPsMzdqcvdXO6yYZtAfhDhwb+JyvlSOCE4b+GgBrM1S5Mep6kW9CJChFnU7
U7a2Hua28osL6L56lXlGthyEIK4NMxsKokkmyaGRhvtTcsbmq2lpuamZUpJkD0Gwcl2LSyexQqn8
8A87Vc3aOmZRL4mCIaAPVS6ADhTSvLJY0kNljsD3FsaXAhAxRSkJupKRC4FQtyuJPgc4cg3L6WoH
KxZqQ681PGkbmXX/d8l7vq5vyOOFOQgO+Tzy8mbqTbVXh2lqEyvDZ/smvSv5fiXdwk+kedl12Bo1
87C4Irfyq9NDB3lv4sYW0eHcAW7+gkGl3VulMH/L1CxbIms5/pw4P3gJaybrN1Glfw9vpSAapqU+
J8Fm8knKtE82ZJh8Mo6KmLdWRXb3LKnIUj7Eex3BE8jIYHKy8dr0de7rrN88dsFWjnnv2eZPWklx
2NCOYGyBIW4EDgOFBL7yjIo9gfi/8LGs3kvnVe+lId7KgRwz2nM4maWGYXSw9iBcEslFNXKo3Yoe
NhuhvN23QDagsgHjbGBP7J5O4ptEYQ/A8o0ZEt/bmKfkn/H2qYkO4ZyGUSeZQiLEv9nM8kaPgswS
e/6LvDkUimxdU55SugAnzisyi1WX1KjStl8w6blhKak39UmkF+r+l3iB4AUEOQosyaASmmAjmSyT
BOFIqoT0PVVVlyxhDJUFaVOMtv++0M3NXJIeOMsVN7gnvoDQ7QjKItdtNPrH1OiuObMe8fQap08N
rzUx5aovoYQG3EV2NAKIwrriJllR/1XPcb3iF264slDnGErTxOO/dfZ0FoASToZlFdW/DBAJtNfA
AEmG/04gP/eiV/SNT6ZEO0fTXDOonvng9buNPNUnvApY3ujNh+OdId0Bw4nA2LYzgaU9VjEqUukl
35DcSw5mN898QY7PdktgXioNFgQcbTHQScDiKwoUo7NkOV29ZudQQCC9JU1WQQQL86xbER1KQLAM
NmEErgTV/Pl2FUQal4fYEH6zRjPlZdByag6xvngNH3cWfUPF5ubDiZnzen4TAnLhIYJIKPC1xQlR
+lJbBVlLUW/JXaleIWRHeu+xQz8z9lt8nj/++0eYJB47eOuXaQyUDhhoTpla+nL366pg0FK/vriJ
l4Qy3Qad5LWQbOuyxs4BVFgQ5dYwUkRBg7dgGfxqoHBVQ9jKQUNQUOl/xP3Gzoz7eJWA0nMb9hk7
+9vVyTp+yPlR0icAty916O+9VLWDQr9Rt9q9EqJo/Lqx/n1OOEcsYmMGZiq0/oXPzbQT1Xs54lQe
r/Ljjr4gyvaYXzm78TO2m93+qqmhDDXaw4xFP6HeIWCtMSBn6yEDCMG2CDWP47kkZ5sS9AXTSPDm
YCsv2dcTHUPDcfiUdj19kfpM3RG9XHWhKMo8t4aHA/DppzIfcUNNrdz4jRA4CXbq8Y1ahJ34L6SP
tZNhQCvGNP+2VkntN4bXPTCba2TxF8rlZqpUwp3oIfhEnYmx6vNmBqm7BoxZENl2X99frvtyh9qU
Tdx1jS/HnFlDcJQXH3kpeq9oEg5V2JidsgZzpGbHQ3n0V/tkSwwwOZ1I6XKExXCVZ8PXGcwJ2FNE
XXj0OZ67pIuvufxf8eXLh20Sw0A1pPMMjHyzt+iIYOmp5HaxJEw6ryRcAY61UvFk2mAoiPVT2/xh
Urkxa60daO3M9wGb7AaXOxXI953zZNYJaxAmPcWyN9+FdM55OOqf6ChM6rpiEhdykusU1L8aElOS
337+r5wecrUeGQyup6P3suoNkeehktx8tnNgxHOVI15OCdSYhTq6Fw0wZPU7H1dhocVvjHK9WdGp
J6zctMmBoBVdZ4Vzkz1JDvceaS6+fKGR129oc8VasY+N5eHi9XNDAtVVPM5PcrJmk/ihy7gVBdo1
gjl2ZMR69+9dTuBxaKpQWdtK69Xq3i/F7s4Y3OTH68cVvhwn+SWG7po8VYiAbYhPSy06SEkZ9Hep
WyC53JH43FEEVLlukTUI3MaGyhcGT7/HQZCFck0W+p4YLeLotDfj8vdGeiAaLVQyqAnsnd3+7MlM
Q7ogGA5OyErNAU+V3HyzsHzz2a9bTgzwHM7U2Ras2WmXKGtMdMe2apAVWbTdD4z7uiwFbZ5waWOu
45bQrBqbP+mR9nnQb6JEHpsfEfiF8EOFE5ul3y9D7vY00fjQQQWWpjZsng+qR23R1L8s/Ppt4oPF
J5qrp/DCUc0CSAYEKYHFkBXGbyMGJ2/v/jg71OJh0AArUIwO5SCjdMhylwjc0Ux4uB4uDYfmceyr
ZD4Ju/THn0k34sNEFy8e1gSCQ8lX8DPW6Hlpkq1Mpasxf6f60xdC3uK+OkhR3rcyaCfFfdqOURA6
IwB1YqE3ruAUw0kltnrnftG0Eo0cZpQMaTvgpKffrIXNH9okPQKvoKwLkMZsc41aufuqcWzHXEXt
M0CrRPHMLLm0LuAwsluBN13i+3xihn+qgnNJbxYNTKLsKxs/Xy+aJ1uhd8Z62ntQxGisI6XbPFEL
PYzPO13ZSBo+z2WUNb+CwLI9T4dCxu3pyVuyz3wlP+aIMwRXzfz1rkZncOSP60AIrnA0+CR5UdXS
J1BFeCJcAhBXKaUmzOWJFavSC/e3IAj5L616gJcSGew/w7FB4ULlU+ICoP5V8nSUo2S3aUX34cHH
xbpvOljDlC1JT1rQctZnglUNZ4qreQ5gEDqkteAwsafg3ocSMCFvf5j4vqN54D2ogR9CrvGMAD6B
9xpasjam5KbuqclAuMQKzbANtYTI1LCcX6vwA4e+QNGCo8dcsCZ3/x1A3HAOJEZkIU/4SkPIybv2
XQIxb6tw8rRspMAqL6mdXmygF1Gmnjqmzv1luK++wtPoZ0sjpNAF6K3zDvUIhZxa/tYnkW8Igdpl
srQCmrFEE3XOnQu27dCs71XJ6xGNFnLgD1rW1D+I94hSR1gxcUqcDtdOz8OFkSjxCHyfaj/10Pxt
0jNrFF4FiyLfHImGQ23BLpSYkIkw/ToZ6kmrMAEhzr3EUzhKFwJxqq6MK3blEwTOnkRLpJd7bvQt
G5F8aUvnDuXhz4uKO5qXzSiiMDOxKuDRdhCfZpb08cTZvMfCwI16DWaDQsQdlEX6jirbzY5y5nd6
s2pnHFgdzA6EPshih+0EOOpjZY52VGW8fc8cGUs6S7MZFJe9yyMio75wbb8V+BIfP0jQXeiRMR2X
gGxWKl1mA+JMm7kTPH8Qsyk4Abtbb6ojSv964VE0tnSj9iHiTYQpwpwnD12JNvfZ41IAK/zeCxB1
MSnF1m6keq+t7/tvQOW+3B/6WLkoDLBJ1kQwGaogHGHXAAqGeEQFQXVDEkWQaenxUtSJNI+WuYeo
rZa7MwuOROpH3fTLrq7GCvQdThKQNVEoSv8oqnw4yNSpVVePKu8ZbIypwV2jTF031wYE+Q3bAgmk
JxjdaiRw6Zj9JTXx73WTqEB/ddjGo9WfgPRqiEn7rdDOR/HbLEaFJmZIPwfe2KPrpyMPH/zLE05O
lh15ApbykI4hju6RnLfv7FUtyA5ex+23Oc8Qk0Hc8Z2F31HUgigNbLHdaUH1mNHBmnVTu0fN8IvR
HUfwcd5/Bu+h7KFg1pYyM7bmhtwz4mr+vyjVJno2ZE5ez/uIXxHuGMIAVYElfZwMytYcdJ+TcA6T
bFqumQY3im9wyJtR6B8asOxHumB6ZFXHWQKsNjBjk5neiZSpYja5x26PrYQsjofyPDr8bUSH/UYJ
U8ndA6TSUJIaXkRVXjVh3DgpdmL+/8r3OR6+SvYyee7KnpO1WbnCq4OsNol2jh9C64fWYk9ZVSfd
ihgsmgdyCeRXxm12hDbdzWaaoublyVxYm+Si5ADmEyGy3Q06nnlVvOvTMpsvkmFuc/kRtJmYEnPp
g3C3TQ9ShVZDZ49uALd/r3pKgwjd4Oe14cbkHyoXKumECVhdx3qB/4Zljf7x+viBwZ1Nt5oNiBsE
AbvZmRQf91iJiUtNEwk2C5lQc8JIGiUz6wSGV96ZryfgurE5CmmO06XznCDdIyMPGc87RtXDSMQZ
Uk1jb06THAB42GPyyxgJoVmZ4uYQgvNsuc/KmcKEtOmoM0WqZWi7Et6lynhtZTIMDHfQj9UFqRwj
4ehhJgB0KJdcoEV0YkvmeZ26jdDX0KeGTeGuJ6zl3amDtNQrtpV16WBAIzwc8TTXJOqQCMAZkd1A
beZqFcoG+A2gQUKnUi3/kDzfQJkLK8SNLQG/Dd/wFsLPVod7Ska/RbnsKvwDKq7l0Vc9daScw99x
TSeOjWncB4UY2SCCJydui6CDiKbLraiWGhLfoxOwDbZT1pZ8X2B+0peszPgwvExP0MlYsS/wK6RM
p2RRkwXShwkwyO2EycdjfYW59moiBfIgW9pWH+pl6ArxfmOCM3GZFc8Mj7P1ihxlMWSoDVB0yWho
dYFjlf/XihoxlpVc+UlLogzpnEhO04qvoBOau//n3nhpI5RRmdW+02D+aywPEyBDZUh7jklrtthb
UTmtr+bqo872VV1kA2/pBVB1HQQAddR7q8YKxdGQK5ekskwoDwtjzbPk4HOik6Zt6xceU7mJZUjj
u46GPe2v9bkyLVx8zAYRLLGlGtH7pizNSXo8Qfr/GDQ5frc+k9zUP0wunQ/M3jbwHYhwZ56cWuf8
PGzAY+qkwYoW681A02+ROY0H/1WHICQDmDiTuP/C/S03V55DFCzzuXn+e70y3p6zmy6nPisi8dU6
g5XZ0Q9Nff/XETL9jb0wqq6Wn5ddxyr3U9NJXfW/2pwgZLQeDr5/7A+Aoxjivfu5LjeTGbdGr9Pu
sTkRQxGTGfs0NF4E940pdUD/HXgavEsjl4WkaSl1ifszZ0B0mYPPb4PMIHkbgPYwSkM7/NmQ4TxJ
EUYR1cVybeXZ0DkzHeDgz5EBsLtBTmuWfxGkb8lonkBLQ+PaNFga9mx/I9v4ConFsF++R6vRlwaq
BcgN6p5wfKKEG83OaCZBzhA8A9N2HQkcn3Hy+koC7Gk2Wj7A+JCVYZm05TeKqa87jukI/HqRhbl1
P+cYeYYoUOnnxz0qY0gZyqdoD4TVA0L//x4os1zXzinwRPCZDuN94CrHLD0FmEM0WuRtgNI30bcu
t4qjWDfeylBrPunreBrLp2cBhuIH4gT+Jw1APUvTPfvU8I4i4aka7ah1bI3n1L2XRP3cAhj7YI3W
bW+LaiIdkZJMAUTtEa4TpmuIynbx4LKQxShefzGTyvEcn4a/EIJjI6/tFUhBkXr2rXi2vu5tvbiM
Bu8P9wtOU3RBbRsRQ++Brm8bCenx0zu3J9sV4+qCMOkjNCJcuquInlwW5rKEOdozACN1W6rWoSfC
O9mW9srgWAseVZiyeZzkXfgX5T5MfkUIVYW/qU3COb26qB6vX5uPJgl1DGTMBxG+DD2XT2Jj5pOr
x3KFDHI1P6PR1XUkI+zgfqNk7eZrzsHSBM8c4q58T6A1DbdBgFwywuoOnbmocD6yqOCi7n99y8FL
c81aqcWdSdGRGp0Hivk8hghC3ULXGzOhnc2CbxPR3fYcPmRbZcSei2gqEQw+MD9H3EAqvK+UIlvF
n1IVEe39Ffa2idR7QeNcExeimTYOuG+KPG3TPqZbj8cRLmkYTMRbgYt6l+WISa/IF8Wv4cywhUK3
T8xNTAuQot89eCeTlK9T/Hhmzd2Qm4waFk8ijSDrGkOm6Zx7JMBKa9HMQYK1iSFGAIySyGAgUBYW
JxalWAIeJHA1LaAZzkHlgrYk3V2AulCn+ATXPB3VkSOP6KaODiP9gv91pAC3bT+S7FbnAQVT6tKp
VFeTMieQWeNUC/PR/frOPKHgc9FrGSJF4RPZvbqKkAVtHQZ13d63DIVvVcKYL6ZnJLo+9cy5ExvQ
mJpZMX4X9dJPsvtdGWjwXvtYyyY0mgGdK/quUtCGR7i8kLRUv3EWnxJo8vteNauRevHHZMjkC7sN
hEOgGSOEC9UBkRUEF3InYijtnYrisy3KB6PveguP+QpgzR1CQNeLf3FilfhkihHhmbXhe4QBb5x3
5CjwfMPz57ZF8Si0HLt8rOq7zxD2OJLV8F1lxPJ5yQTcb2WR0SZj0bjw8B9s83X5axHoskOdn6Cy
sAb6BfQeYw3gXKjEHTtgG+HNNMkcMAIXveooKXhCnClJL+PfIGOKnMvS7KQkCnLDr057JQjKYBwb
G0hk4nWuyne5F8YVtuh7HW4sKi3d61Jz1nW0Vsd6zhWbbxFy1KvP1vaiNjs8pCb1LOv/Rsb5C9RA
U2rFS9fFhNNkOvhE0D8j+H7PoepZ5Qqxd1o1SFi+3pE=
`protect end_protected
