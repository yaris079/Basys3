`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TS85+Sk+Li+PHAOw1rCfNmgDRVKOnC+41eHBC1BA87hayrIXC1wmU4SvBapP9qpYKhwHwhIpMaZu
js91Kjepcw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E6f+K7VKnxaNdr89s60MI467P3egItQgxmCW0S9T+9acTdK1g0AAhKvSZA/K2Mq0wY6hbYOV5Gk5
TWiLipE21/hj4GMna2U8L7OKejYpiIy+rBmLk8gtKMGOf4k16foYOo+SsyEB0R4njtWY8ryMJPAV
3942MIKZXzx82biK4IQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
NhxWDVwzBFIEmjpW0LAX3HcQpP3cuKe+bKc19w3+8TfCYxuMtdOXO7we700zLbVyIHT2n0GWkJS2
cmJFpIY3Zh4yk55GBVX22YbgUyrSb6DkngdVkFNZTiRJ325owO3deTsr/KtNiU9S7UYN8CewTpII
sO9mmEC4jZKceDYD3utH51Ga9rwt2HKYsT8LrEb2Xoxo2E384TkaLAaCWwdaYDKMXCrQwhqO7ZgH
GKXA79bsIEijcjr5McC9EZE2OVYy3oqwTnbpF766YEreMk7CC0hZmazFENAS7YAZIHn+e7CjUT5y
h6B4vr+NKDa8xjMivVgoHQ8o1ulJm/5OuAB6vA==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
zs/COoZ8xYohtGibLjBNGCDTij5Xbi2eCEr4EWttznq9L7kCO6Qv+GSlj0JhRRSEiSIcUPCUPvSF
FNUOmhVGY5rCEBWW5gPs2U8261sujX3IcKo/JPsX2RoP2+smTyZOvdr40nXpXJAjtG4YVCIVPKpb
OMuSTjOrEeoG3PtyWAU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jwZ3f+Z9zVxKBms6N4dfKYbsAYphISuHtO8S1nMEMdL3C3h6aDZ1a4GiDtg92a+JHS08kN0MvRew
20Tk0BrC8f6w79fAhxQOI+DmOKb3FB0FJJB1eJRYpVI1sPah5wH0IRPdL1/TDNOcJKyhWZNUjLdZ
o1HexrUHq3+behnsvhYEaMWXVrAtF4kmW0m7pbmya8+2M2oOtcs6gYOy+FD032UjgvMeSvYdtRUu
GVvC3V0TwIYeBz8tEbJ9lNJ1h+OOlgguI4CbuuSqbm77gHcg8FA3G/mlBYTHIg5MjZASq6Qrq6e7
TSlVYH49iAUNPQ/AXzjQFe6+nY1YZzDuwsVL2w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5200)
`protect data_block
TC1iHvNehHCY37HPHPEf6dvFlXLWF9D238DdJ9ppL9z/nXIo/tUWvCgCf9PtspDMb07NM090SInn
p2ZKIYfITUELwGKJxDIlJdAQQpWCQg6mxkSu+3oxlNUS7V7E0kLAbh92H9h9Pl0AOB6TpGyeNoka
74c5aECGZGR5wGhQGFJMtprlXr5Vv6B4pPn3UTN61N6Juik2cwpgZTCCf+TprbTXpbAi9kz0ByhB
JiksKBVrjtBiUsmdif1vhljACpN3qY4k57UPK/WltVjQhAE9zzfezgB3Hb/DoGwJernAziC0/1p9
upJlbDI7yPLIMhqVyF9hNdHc95y5eyvlbBfmkd+6T4TM+T/eZkHzLQ7rFypcZxkhrkmjSc9cvAky
sIdAnO3NldGpuwbPLdPz5kVgl0QypOUmBmUk+ZBN/HYhLhMPSb7uFhNB61rdelI45EOcOGThUn7e
SL3gE3YXW0/jU1XOOYn2fekzsnsTGIzOMbAOmsDwkxeF1u8BMyASKeTHOilkM14Yssge/YU3cflW
PGrKSDmOKbaap02xHgED1XVKg3buVpODOghP756i4BotZBgBLMT9G2l2V/SwazWtGOHRofplQnov
rXhMut+5QluJZbMA9SbfoClPMsy9KjMGGwP/UIZFCboP4JA38m2NC1FrW4kmmYeyhe5N/F4Vhy4j
9qvF3brDHkVNREx29OjoluOrc6x+JII9WHXdJOBUoRlvt4e53Je+pQ2QqvwHJH3UFD77NSLXT44I
s5orC2zZz0vk7C0sHjvgEmVf0YRsetMy7O1/4x7+QDSoR6x9WFvz0vPaRT5dXqUZsG81y2wGsJ4O
RTTlleLdqEcOiYhVTPxkyU9b9YS/9wX58UVb+AVH4ykhWfRgO2e1IubbjkqijCrCG6OrNK8s6jUw
U3+WRid2Z2NbcOTBX48pV8I5QFMGi9wvK9VKoP8diIutORBurEL9FS8CKHXx7bMM8CPcPqstELcL
Arpi6zUTseQ0CDTeNnCtRkgfGnH8/zcZ6hixUWtItuh89/9i+p9CONzEAEIY5JTRgPsJ5E5iQKVm
1sZYFtzMwnW59WyMY0oz9Xpk0MmprA/1nB9QYk2rZpUGgSJC0LbRookfl0+RqG5VjtnxGerJkSUu
BBHXCyNMvH+gSxrqY5kqQAfcsqzhHqndWYiPzFjs9skFEQCOSykLxWBToSu3JqVQW6i+d+L9hQ1R
gsJBjTe1Pvk6GKHP3KRwd4ZeVvttVq3qKsuyQ3+j9I83Oah2wAKjabrjeCE183tl2JKt/kNQ5Do5
DJSSxPlNPJuh/+HZnB9l0k+1HxG9eq9KJPnRTeDe2rP3obaqFxR1RpbZKe04hVIiae3cXEmC0mNg
96cwsr1wqmSeINLgpVyg4xrTua4cEyaz1TBlUoWXeV6ASFfAE3UpnoOHqybP30pAzYLNUebQGyX2
970j6C2ot0/yrKQpDzF6HmQ29IHWM+5oG/50btbtP+DUVLC8kpcQoiqXXiV1eIGwpEun4ccLEN2s
EID4xueTKQGUCEeNiJ3+gilqbU7geyqTEgt/L45QUIWPNoHDh15pxo60w3tCFQ4Nq5N6AwiESwM7
uVg0ZxD0z69X+hoOJAusWZb3sB4gUNvHNZbrA1zHVUHwkaFjp3mUClZlBPk3fuuXWhfZk3YjrSpP
lavxaDz1UH+x0vjmkTmNoLvOZ1+BComcyAk4fDuGgW3o0mLjrrqmjF0dwMO+2dlk8AdVr9ttgdEy
l512SJIw/e7ApV49X4ZVqOkRi+xR+OmBUbIyF6xCJLF4kOMiEU/X74cctLeWmAIAe2HLxM1uPrhn
Fy0al6SyCV99Asf6WiZ4zh/0i1YzLzA4YJpnW0EnnfHTmWUPP4zlRIHC8FU1AlMZ1Zm9rQrXUwup
PUjpk8j9JOsarG+U9uYGEh/VH9CcTFijrN/2tdyRQZ90EJhrDcz83j6ZTbaSyiw3KU3MnmA/AJOA
hUedCm9z3vYb4mK+pLNNNcDtBSQJsQ8onb/6hzRz013hGiam4x0PKIl3aoBF4e/P+fuKVueucCLP
XCHdFyyNK3jIYK6ViFAiqTTe2N30RuoyMTXMb8vUEv1uI2JuHgQb9bUp3iRNcPD//uTmReHuAYwR
ZYsrWQgdJufFSz3jrIVPVu6K0fKJ6bI9zfHsWWaX69cFlDl60L06lknOTAYZHoG2wQ7OKl1EEkIn
XzfqnWYG54ji38kOp+RFgsyXwH3HlmvMrfeP0Y5jf2/0OCZtZWcYVA9nxJzx1m2qPU4GCk7FMVfN
hp+BtEG3EAVE9/Z+yuyPzI3LUjMp0f6wZN9eZfcVsQEFpG5wm9prFYqYi4nxhyCkxZpG2I5WWMs+
iNPJD/AW+ev5ZhdIKqH4Tq2TyRt2Q1jvYtq8S7wfhSZ7K6Lx+13CHllf/PNPsSqVrNwDtK0LtHn3
Wc8OUGc6p1sJl4FMSCiMQd0W5Cu1gBlL5Ba6yi/2OQpnyt3UHKsFBdksbDUnMN+eQx871IL8AQeG
j/bl8YqjpyrUR57aOK2gTYp21vKa6orS+O8kQPu+6DltTTotd6aPvqXjnEgg6Rntf7S2iCOr+tcX
ZIk05auJUcjmZ9SYF5Sr5XC0Kyqnty36FGGQfNYT9Q0dtQeN9gpfojJHHMjtYuGkUNe2i7fXZEce
m6PklzTALgCSU1fC5WJORg45YjHIhHIPEiuU62eWLiCmZ3L0d1TlCPExkLbLZGRx0fwEM/DSTRV5
4bjPQuWXHQQS6TcGSfhUUYtb21YRJJ/edwogDxgp6kYHx7NoOjVTCzlh1Dzud7ebhimMa+HxtLSK
4bs/IWXEetMInHS5WY/MaMafnXiOJEQwMNyMZS0w2oD/QNdKotIO+fhfKQprFTNGRHBgr7oxJp2a
Wf4ib+a2F/2taT9tb/b1YZ+8BFGiveYFaPXo8qUAqhhgOpqaaSyIGUkSG51Y6ZwKF3fA7BZlr3+M
TG6QmS1mb0b+Bm+kyBHfINpg3iHMvRvm8PedNKfYYXlVRWjZkDTn8kcJJ8mgQjWmG0PgVbdpyugf
qQM0RSdofivBwbcNUav7g+2zA78iv2NHPJqxrHTQozoo/a3/VoRboHCR/J5vCN9xJVk7gZ9vt6Ex
CNyMcQ+QUrwT8n77TzMF7EcNKhnGkBZkMJ3+6wi3dR//oBVcl5mjSvF6dRUFdpHfua4TykRg1amk
DpoBAQRP0u6abt7jCmeOjdr46eYZzIkK0UXSCLpM4M12HY4bkw39sOX2+QGavWQza3RVCIBumBXm
md8gPhCPNvplYIEYyf8fR1UXTYvsj4TMUbKRqH4hwsWfhU2/9OZ+wF3/wxaE7mf93UqIRwS5mULy
S2qoJMJVuHpRW5057xzleuIui9yGPaOONkLtj2gJFP9Q+Jdc9RrcqsvQe9L/jGY84xMVSa3LAzLt
vVJcEQDzlOKx1pYRdljAis8wbTM3YSdG0AVFHLeJCSj/0fxeJXhi09LCLNcNNTIDfjHSTO22CkgQ
2zPbZKfrmLCcJCkwg8IErKv0ApkdzUW/YFS/d6jd664oncCdFkYZmAn9ZZi3QoNMoqQ0T8Iq/GyY
VgwOTKcjEintpLyFimtf4cyF1Cz+YThY/fO65GGtHR2X5A6nOIqYJSaskxg3Pu6grCLQntYw7tOE
9ehLN4GYnj3qUI0VxRY4V4k5gQYFjgKpC3g43KdWznr7Dnonb+iS2MPhhavlMOxsaw5H4PUt1Ra7
tGP2CMKZr4PHAb+GGSYf2OZgpFMsrFU5COF3jKFNrHGfxQgySBl50inZu/n5qmi9Vnrbr4WVGbmR
ubwM3r23+/+lahvymYXuZs6unqOHlogx260Xe0O4WwpsysRrhwXNs1t3jJqNdSATOsWgLehoJSVk
vB5SvwddrYxxOP4+D7++9kgI4ZDEYj2UEuJhMiR5XvoTgYa9sJLeznmZcxRAsNjkqD6VPNVv22V4
pNsc1SwSHnFUCGv0xouAb1+q1nHbo5jJ8hteQgwhT/eXdv6XNKjZYCNDZIu11SIXj/XOXKfmPG/W
Hf49y+G5EJHiA/BBc6hGWia1Hp0ip6WXAsNK5AOgNt5imZDWfPQ4jmAwF7QcW1LcIvKvYv+HW2Ym
ptNN8x8fQH/AdtGkaXHzoAF7KmUvaEnBJxufZrXEu+MnURMio8wCMPKz0Uzqjdu2pNeY3TFdyQyf
W6VmiWuijgbciyuG8WSUggLrUEDE1MLS8/LyEvlBfvztrbIEYrIDkegHxtXlXEM1Ta7LtG2pvJCa
MrhNS7qg4HRdZcPgyFL3SYkJavrkd8/O/BZe38Hkq0kZO9z+9gJpG4zY/DQTpO95+jkWHPi66U4U
+Mq8qajz4UaRcoo9PGjM4qworQXTii2W6DKQtCaGd0rPpOSaXA5T5PDE4IoRfQUmOrwLUrFbv9Yv
rB6+i0jvw90M9oSTsQ3mWiD9f8CQBWcS0lQL9QRDmZ7bNjeityTY9T9NfCnHjHF1ObkK1/txLUlA
DQQ/fJ9LDkeIwTvA7xKWAtdkDjtLqCqezQq8Tr2MJqFFiOq52TFYxam4M2ciwbSxDZ1P297xDMc1
EPckhLsu6KtpVc1Y4gZGd9EQg3E90jwxPC9S0KVlIukdRzWpU7YNgMgYMKbSNEz+hBU+T1ff8xOy
wSvM3oEXEaAid9FzUYXBU7nGshhmjGzuDGpiyDxfcoHK5UdKjzeabi/NkQK4DfWEM/zj7VkBjJVC
zbhhpyLtXvLzmWnCWOLoQ+YJWPWjJTbCwcE24vAfbXJB9RVMEF9UAqIoLo62gJKT4Qk24uHt5o7b
2MdZg3V70keh2LUm3DahE+yce6tkxATah0MPr8TQ/CDCiGCGH2AE6GG1fOVpYAAgXdLyEEmJkpD4
2wCkocDg/l4S46XuYtOhjAHbeZmluG0+sQQUdZn9eIWp8UOC67xvzzaWFXuNoJZBEg+XftIveaWn
isnIakprXxSMfssbVzwLMSOlByGPSI20eqnh0uz6TxXS/NAxqz5twtLUb7pjraU2DABgQ3qT7OLX
FW8F4+3gjDUdSw0TMJ3BApsmSku1VmhIzCKpkYdONyjZeCs/kk7byp+ApKOmm5CDeqZp1nqfapQL
6xP52sgPDDlThzZKlL26RsF4GseQe+uqFQam0uzS1ZfBChNVacgJuXkX0jKpMpyOgfawfSI54NHt
DMf0BThbXtGBVLzIuz8V64ECCwZ0Ix0HnrdycpVRhkwKwnVzBydVH40vLx9aYwGU/39bkjHNh7Ou
TCOILfkMkOPLZY4PFTuJ3WVEucvQohz2PkSxPszrafrAurX7wmmAP6YDrx3rY56y/7hSpHIMn8IJ
a7e389ej9jUsEbuCnELAcvV5t94a+/MZGJw0Nt3Zeqx+uZMgagvtZiebokg+Un67r+nyAdnhnveq
w007X5oe6TGtPvBUTAKSL4Tg4YB0VtL/GXMJ4VdOXVvfWK7vWi+KJ47pxjkVDd57WYPSSNFZZWaT
cAxUR5EWX8gVLCbn10EJ5j0ZZuyiRnqAlFPr4nPtrKQTQpZsf29lVNI1iu/tCyrxhfblWipPseSh
fBi5mgv1Qn57I7sCSCvsaAlpmYDl5nMjhgbxacm+EkWC6Rj1oLQhK8k6qACkeYOIwUxZ1SOVnWeA
Ho5s5JKrbielg3VwcPfYRCGfVWnzYCGfTxUgw0j93HtBN9314m0XENU7lzIZHe0pXbmnTN/Zp93p
4Z5qZHAsz3jJWk9CVRqqWFrfuE8JgsIcubO2O024YE46/vP74BzjlmquylBsdh/M+k0NyQ9PEA1W
iwIcS2YmBpZRU3HrrLEIEPPHlDfdoioT8XapM1it9/hN8rB4wsLs8b/rMGdMOr0emg9Glh1QxqIp
S8feNYahmrZCLcK/cnrZfmo9VlF4xZVE4tpxsTdFXABRPRX6HpPQHkG/jicRcGn8mdGvu+hSoiQS
B6ubFYMpXPI2yaPUpFetWtGzCQGSjq92sHBV77M+dzxEY4vQhla8Rki45i2t3RRSBvHUN8WSic9s
BBf7KufIUoVNxLccNXmJLIyaXR0+lUzVaZkfjEPrJNVgD7XzfOpaefdILFEI2MHUyq32vfesV/X1
DAgfgc+j+vggM7YDWCET9sn/2M+JcfyeYGx1/hQAp+y+YuReJxRVZVCqvYPBw09ULIbBpbp9jjgz
PvQashpE4fCmCtWAXFwjc4PCCvaE3bRzbGOgnG3mFkE3EnjI4RAe7uLXuVPCEC4O4fBZaVsgNhaz
10G+NzQd1drTrxseL2lOROfwQK02hLUNHfG6Dbb+MXHwDdCBaBuAn7zTy2YqRRxDZFTuLCc+mnfh
pfbhbP2FxpUX+sRhQzyBk5rh1nJqLpwJFLK8av3LNV0lSFLBR5JpYPNmf04dkoPyGWUsYFkDPxb4
3KnFZpGJ8ibz0qBJ4DwbDQ+azJPJd6QLpfezZv7sxD3PbLsT71NL7RfIyuy5vtBICCrNe6uL3mGV
WQhIR5pDpBdnIBffKmCJj6+f1IazcKPNFPOEela2TrgQYKqd64NFM/xYLt5hI4tektDGxneXrbRZ
1+G4fTpqJ11cKOn1EB7+mbxDNU/wKQjwzmQNVhaSV4F3kTwmmsZU/5jrqESSRiI13zC6Pza5akw8
bEHHg5nmyPrUFd85MtMc8PjMAEdCRxLaBdWYqEFDxAkutseVtlYcW0wKjcrziRBbGbzvRKpwNuQ6
AzYrQFmktPdf9+VrUQvWXALr/KTOQ7mR7+3pgeUEC5zIzSYFkVhS8zNS8v1J9kWPwrDKnN8alI9w
EtIagvO5XbHc7WUm0aJx+Mf/4YkGxWcev50stqiNu1UV7vJM5776dUil2sOaNaFuOgDrLkxogoZU
XWl0slq9oz1okQo7YMZ16MZvPXD7gWadLoetSmGw95UNM3RnxTi9+uq/7lE0wWsTXgzeSvQpT3k7
w/u+oNr91K10xDAKUw==
`protect end_protected
