`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
N7kVdrf2DDc79E35x7O0uUC/PhkMDVIm0Crphl2+C8VzH0DVoHa4h0xfOLEgWX0X40HOcLqHYCk+
zhcWlhGhJA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
P1kMFrYg/qzqMqCMW8zBdqd6INzyGTJJ3mS/5p4iio2At8nO14yHSvQjs380hxXUHs2esVK7roqy
5T0xN+Rv7iqZ59E2mJqEbHyNnbBlRF8bvJH8uSk12MbS0vlbc8m0pCFGZEZFrJdIJin+D9mCo/h1
gTygF9aNngZzXI84ILU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QlUarLjPwO6swXxWGWAHQ2OKXimxp1XIFh4+fJhtZGhoIYxmV1k8exC35tt3tbY0lnQdRjtsOmT2
jz2uEycewx26wkNPY8npwS4kYw0+a7GcDPlxn3ojOw5tr/MBk8h+j5WEN5JKXd3Rq6OUB6vwrgFG
MTNktOtxug31kLgQaOWACLVUvSd988MiyiCVwbQJ2evpS+ZM8eYbsKx1+lkuPbhPqE1Fflpp51Ht
DXiITvIgLAnkBNgJnyYLI1maxA12EzNDugP5jnt6+pQxp3NjTdA0u5sMVZbBI0UGUOQRFJ3csuCr
E/kQqUO4iEa8N56Wa90TzHe77wTqsNZJBTuBNg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
f6Smr5FYSbcUAGnTEDHmFSQGXhB6xnLo0/fwHOG2aQz309fo2CJgFmOyVagU55aLufQ3UNXf0ZzL
PAHA63YUA5x06hJjV7Q3OD9wIdBYL6541Mcg67CHYBQYU92AxsXLrJpbeE9Me3u8XpPK/2wBANRM
ALJyHUB9N0d7WdtmrPU=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
sHoBxxk1ECxq8hNKHNYZ+Y9yB7+ncq11V56JdjDib0BkEATSM28xAXC/AzcWI0plWIBzPb5z15eD
c1aFPGsvFE1heTxsJMnqn8TqhwRRWbYQJlarg46V35EJb1kZze8/j+Va0UJSAZE2nBfNcp+ADRmR
KSyyaUrBYp9VbAXrKpcf2eolAGcnWc/+NZ/0voq4Z1nsg9fFZ0jNHGy5TOR8g22wzCp3OF5CSfK0
4WkUBMJqxjZy99m1arM5OQPuwtMh8wfUn4ez/Es3DszxDVlLgDluTOK8dsx3E6wnhrEyVTylXiXf
3xMY4WsWRZn94CjBLcpXHGKrBDayGL+uIzVwPg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5376)
`protect data_block
bZTwgiJA9YPD2+2fTDNVAr2UCOLnT8EaWT4w3GQX6NGl2+4SpSAeRbDQ9TRDvah2n+yjs5jBXLXX
eJPy9xjzWTl9ImmOiCmP1fFEFHCLZl/uU4A9tMEM1EDBRF46Nw4H7riEspoRT0PUVGuS8oKXzI+v
Rk41yYdd7p/ZavVPFQ/9tNzSp3dOkgdPCfl1XFrYxnjw9c+NEpWuWo86HGYILANVGLzlh2aWh1Yt
pFPE5woRD8cGF2RP//4m4y60PDaFEx0tKnWvz3pGyuJxkc/LDYXrxavYXhHAMqcEZg3Zk8PcA62w
2+pf6ojpTSrMLWizqVCmbgWtGoVpF/EbTEk2Fv3zBhmObd7yM9/j/TwQAEpt/cWi7GieL8jZnh/6
qJAXRdlg+eRfB+lq+S5peZBcVwTwoAb1aAziZG5Y73loMabJlWPS/624KfSWDqXrFnrJWmOqXBPo
iCSEQqdO0nq83ubCqcy7YsZMCY1ggrTJApmLRNkWJSmnI6/GwYo+yQJ2rKwKvoPnrdywLpVNruTF
XR4hVs6kQBji9j8zQebRD6rxF40d8Orib7WxjEUwgTSTpLRu5GIoCFU+PTks8GVlq2FIzKdqsJZT
j0n4oVOewLoNwm8uqVz//r4Niag6m7X3D0ibj7tENkh9FKkV3D/nYzNVle/dRv3ME1V4osQFTqZ6
qTSTZ/sYx6Jy71xtAVxSW0v0feRIms1RHGb3x02eHr492Ib+2S1V2uY+Muwwt6fswQUN0ohCktVn
9afh4FR85k8GmKmghxXR9bMXq47XhFEqZytj4yMQLYzPTs8oKBiXPMoiXHnitOX7Jj5df5iFeoom
wattAmItzQVRUKYGxY/26KDit6Y9VK6ZD3JBTU/RNFVMgpHF4X+SYrd0ToT2NeyofPIIfE3X8Phr
nevI5FSK3qlnHYPHBd1tsBkyhE5wfErvw/LswNW0nKz1o4jhPj+HeRXAf9ixbBRa3LyyrJTvt+BY
gZPRE2tCbB53Oyq49zajVmv+ahXu+gvUdSSmpMXkecPW27CcTvFSB1DJgVBQNCCEV7tg/j4jpLgJ
6YtBytRZhMnBf/Gc1GkyKjPjARncTKcw88fx/JgAxAGDEyKeHeJEMk1AoSAiSJMogV0YxijMJU3q
R6sjCtszz3CV5k475Nr1WYW6EQP25m49C+GqvKlmnJ8MISuotpcc75k7OLaGS7KCCyxSI0MO7WFf
8sj6xmdozfOv9L1ELtKYxyP2rKK1NexvEhsy4ogqBGfgfNx4FhjRTTZqb1Ma+uR4rdK7rg1PFkwL
W/8bvKgqcoJoz1IJoO+lI6R6c1tpjQkSVCJY84GZ5dqtjt8J3QRMjKwYOYczGALChX4L/bciZx0h
g/bzPxDF4lr9RP1yhNE3r8qqQX7yM5zs7aONHhnhd2dhUlzmekV4ADxNJyWwXzRipxFkIRQ6Djr3
Mkzie34UfT+P8rS0+K5y68ymsf1Ldg4m/RUrpLzwSjSI3zGkTJsarOzHGx+zZLSKYSjAK2VFYGOv
QGNRpGNMSA5UK4LAdVa2vuXj4aliZxDnWIihD3sXXkW3wH4ue0ZPxcK4iwgEXXzgStBAFy012Cdg
VY86uiwcLhMyiEDJXXYdlzWAeU6WVwVVS+vXW2QJR3ZXRaXTxsXWXXBZI80xU0/L4HlXRdgMq7Pd
LwISkZticDDEX9KmM4DPVhSNMrkUw1x8hsruFFPHxNeoujNnXX1Pt6KYL6rz7rwQufKbI0peygyl
JcuQmnBhXNZv5rJY60h6m5cDMjOoA6hAUScQl2WSTht1CcAo82iKr4K2GjNL2mpxP+O5Bes3TeWW
EXN4j35fpwvJX1imrJ1Mwbp8o6p8ZiN+Yhj8RxX6kq/PuvaM/4UdRHeyCfWemam1gNN3af9EIAb2
YmiuuaumfDSLbTpbZDt3hvg2MKIzG7O1FjffbQXdqlrCSmYI3pVfD9NgdW03oHL8H5dzLYSTCnj/
sWVERe9ofuDO4LsIPJceqE2IjrRCdarljqL/izzHqO3p+DlhFTIgUP+DI27JDcT/c4dWOKGZZS/i
hlNc40fo4NhZZ/t3tgcLmysNa+llBIIYhappy3xN/Qncg4Td1ZOOakX4oz9vm5v/B4A5N2Ma+Pe+
tAoXje7y4d/A3hw42zIUbKqhPud1KOlPuwCj7dqO9P3U7wFOwL0xbzmIqJc/bMPcXREZik5o1Rw4
uvLKBlk7aUJ4vv8xU4jSJfTFlqsHgUY8LaKxenJBDlkbqmHO48wUGxnG/zFTOILHWj6zIqt2G54+
Rr09xY/F7YmsDiiu6IjCfGXAK1/003xW3jcJLTyl+qUFOdSeG5TttMt2/RedjBeZcGH6iIILRG5f
0RsybYXqzh+YEvVhKZDMx7j/63HPbQ+SXr2TlrJMvcjw47q57u5yZO+r7GEwvILf3xq9jO7g/G9L
QgxMJnWJrBkLFezAGSJuu5imZ8v0aD3wicczrFm5jBXVkXEVYN2IE66YiK6+wHdTPOwuximQHKe3
DAoZLDB2apCZ0OA7gKgTF9hDYY0QNQ3m3pa0lI0pOHJMULOqr4pGlIaC4M88SbcENnjDCSTuRZ18
REle8s4cgnJ5/2k4zJOq1i3tpcSebMqnWv30zwxgVf/wXMjAUpXBQXn2I2zNffuPIQPaA4lZHUaA
2LAUa4LLSua3+ff8x2YwV+T3bpJwFsbip3uV0L8Nrf21Ufwr4ebxn6nZV68Lf8cEMkJOx00hc+gi
JICgjCXqdPUGHa7MwXT96FdBIGIe1Dj6eTFr0oVtSLUDiLNeji02yxIguD9cvfxhoQXp+It89Lsh
mW+7hMybaKfm5UNJAS+m8vW/jkrU+QCwHtEaeTVJcVxmtZAF1JujuLrhXCJUwFo+49pdXhj6mxR9
PLhVPRleJeZ4lqo6e4ADDBJ3iNtznxsji89+fQRi7flOLAGves9wsCL3jwgkwgTH1MPRu0vIkMjd
FN+8gAVoOkc+1cXSCHY3X65WaP1nIH/Q4nELw02f2p222BsKnn1TwSnGpCRyf+hO9q+HjWWhx1IQ
2pnqnEFkIJwY7DymYKdaJwOeI9+w2JZ8vbNRA6xm1bqBiwIjXUCxFt4xesaewM9lOaYrGMoa/pLA
nSLDZxrOxstr6mr9BNt9V4An+LT6SoJtWQxPBwqY2U0C1X03uZo8ItcOMe+0Qy6DecswOfpYqdrN
YCKzPGamo+frJvRoUkswl3E2jUmS4qIue9Ij3+SUsk1Nz6+XfU/2mFgfr17H+DKYvrYNq5zkZZ3S
3+l+HkBJpmirf7YYMa0s3fPNrc/4glZlbZEzVfCHcrQqSa+lMl2+JuDQ+IlM4LRzDqRP9g7hq6If
Bpy6+i1g70uaWINITO3dBOnqRRNmaMnPBHmiDUg+/xm8z2O+Jm1SQqo8b1p1bsMukkryM5wJiI1a
xfLHSqaXRJQntcbv9uSFtZTJqGhzWpQxv9/HCn0lLXjrzcVOXSrYNciJssTEN8gF8wZha58z7/Qo
E+1YVoHjGu5Do1LDuKryG0eYt4pthz6GAKdLgE5s9pVbi4xfnFoX89bOmdcHzs5upg6zfquZJjXO
Wrr5CkpeUySXJ7IHYK0XUsCaCrBrt7sAbB9IWYBGe1Q7dg+N9au2A74v+wnby8hdhI5eH7YPL79E
jL9Mv2RBmhb/WM8Sb+ht7df/11R0RBC13x1+0PB8weVlfzJzP0jR6QHQ+fQm+WqKWPnDHldOj1WH
8nYa+TLn+L1XmXDn3tYXGaZD7YeBeodzCcDP9rDXBZn/LOWB3YkDSveJVdjU0rZv2YEbnw9OaQB4
oTxaF0xMLYCAnU83E9gkdhQy5LvaSDNcC4HrzAadpSBVS//yZJ6R9ZIIuf7NGFF19miEP7Fe2X3Q
SW9ZVOrSSC8s+3NqFY811flrIVbNfTSWzTlRMXTQeTPaiY9mruVzc5K7laG4oM4LrtHODWAX2EVS
14r5N0o/xM6LjiqV3sL1acDMm7/cO8KSq5Aor5immsfgJtmesflcGIHpXoASQeLAwrSu1wakJbZh
QTyT4ewl5tHUH4GlnXzyWG1tU8qgl4WvNHsY5djixvG3ySh+GLXwMtj+mDnqLrw6zryTBQb7H6kR
V01b5qoTMCsdeZAjafZOPZa3o3cxjzn6uYlNEr/UPwfy8PPM6rGh6OgYRxFmugODnwILsubhSNDV
oE/GwvDO0qNUAQD6//H/+F3CMzUGj6LDLSgm+z6YVKb++rE7Nl1RM49rYSWWSIgynsCQGwWe3t3Z
L5Jj3YqesziN3cwaF1JUzT4fZwDK32ioaUEr97oFe/WoqDWvg1YFGosH7Gy2uB/dLEf1nCi72IiF
iiNosuQdsWAcSFNsD5vGkwr/JVMtSYbh6ED0k3TwKebBJ7TQMc4W4Vx7+ZGNdlOmbPFVxQ8BhuCs
kTb3TdYym14HPTmZHK5vRk1+ejDuMJOEUIxXKkdnfxJxCnRWhDDGwYj6Xbjoi7GXsVwq8MSl0YCv
VeVo+Y3uLSsUCtHCLDhdP7d372udYDCqa/2HsWONsaMmPMV7jaDEZgERyjRRI9XSRXaJvjtOHINV
omL6+63BBjPim9rkSCymDR/BIUbOKd0IOz35MgD2d2p/LPKmIDrR6ar3Qf3oFaFaNvQDf8Kj7Z6y
wuG2pjmtLurWanVwXmBjWp/6YIla9uwqyjZEzCNtWpd5Si/d0zR2I/EOU3I48bBYo2WGZl4PHRS5
/WCTc/QII30gmQfvcF+GlvF2IUzZL6rYsFfVDW2GaeK9GrSSN6FRbYy1DVZ8SM7tD5BaLeHubzCq
USU4gSbRpdHC6HNipobdBxzx+5SZuEa+vvWMBpwkBLU3v35HOIE5hsrUyqbNeMWuNbKgGEsSGnL8
5rrcmh+R2vCyLaETeMYR1iOBbmGT9xWdx5Lb8PgZ3yTKc2o5BmZ6jY9WZ5NFKFNvx/NjQaKDmV7e
aqPjDvfof6egahinFS2w3erWIjGZfez9uBT3E5RtWTJh+4n3ZSHEvniM4jod7GkBki2wc+defZbM
1+lcIwSNQlXk4c5yd+NOGaRT9hs4kZ2ncoIvPUdmbkXYDhFhPhf/+BJBAXWUr0yv5XvfztRce+Yv
4RceGAmPWHKCPp7wzW+CMXsNcRtnaGJuyM4ijkILnztNvtfAF1omMtGKPiyRjtpZqQgfN9b70Na9
XnY5vplSEeUnmJL++IlqOD5rMirffUDJ0pMMCYmgajry38E8+R+NmrXgXXBNw/LyAXsnqLsNq/Ww
OwdXuSZnlDlSOpAlzNhgthBn7Nq0MxxFhTd6Co1I7XpazvDw39kR+HO+e752I7NYiER3WRbvA4BK
pzASVCfpF35UYU6dPYfoKfU7g4sxARlTO/xevgJOvzlivouUmP3ypojXxDZqXvyul2DyEn9mJqex
sFmgH5ynjCBpWimGg2l48zh47xnwa5nlRBGAHb0gzcvRY8b2M3BMDXJCkIXlgYBhVdt0SbLpmJ4w
Cts9d/D5twLMfHti2GpC6uuus+pMKvWp49f6IdwhdQnMQqqc5v0IL3taq9cOb/X8CEoJPKVJJQ1P
1N1YDGEqL2N95PXj/5RCo4mJINUqtskWtARHOdR90+g8ZArxNUmHHOrYa/ef/3h8QK579Yoi96JX
QfJEb3wU+zOpO7TD/4RQq6UscMBDQHJXWPI1wq25Yr+XLxjJhsENn7LQGiBWr4iiQpvweHOi/ANf
+MKavuI+2MbCzkO5py1bfsH+IN6rBs7jU7xKFcW03jWrJpaLEfvIZ0ejHSmFUyypu5qSZUeKbnl2
oiFutqR6QEejMPTsJzcWR+4uL4NwozVPAPhJm5kGxjawTWqCxYBS2rEtFxmBpdLudp2IVGrPsxsa
HXDdB5e4YRIYRNma0SpTK5vz8gIPgp2AP/5WPnn3u1UPK8kr3s8iHY73b9pqzF1qGUzqIHllc9hP
BSZivf+V1/qHoHkvsqr1nYQj2vXimdcPVnZpFNbOW0I03DaAlCDYhKwWH3Ru2qtyrk7+o1oVg+Ig
QwMuL+8lx6cmpR/62DODLlukacAizKEkEDiw6G3zK9EHwd7Cwly25gAn8nISALvovxNRvyzdipAb
0cNvM39xuwwDQT+1+8XrzHrpKKaxKi3RZ8EQLYfOwRyqkHNdQ5sc+f1WsV6WS9hSq+9h9Oj97bYR
yfHmD3RaXCu51r3Y3zv00OWLFLWn2SXJNbQBklNzm+9yBkaktplGZ2kd+kmUzc4cyAl4DEayQ4sE
gy81RoMX5Y9oTN/mvBs+Z7TwutejJQXhbaoU7WUxyN/epKsS0iK/Dg64r9K1C1rGbGhqCdf0sa9l
AToCU8pyg34qllVXm1hQ5aHeV6GTL0LimOlPUAdXiVymUPr9lSHVyutGTJ7PEn+YRqIARRCVvbaF
YW8Z5fCBFQh7H1s9Vv05d4DqsYkJ46ZErifnvE7pqbRIK1SZVP8s+Zz2ShjbfymzmFW62PtP9j+5
W7GFDOHBXl3OKUbHkIdKP2R9tWE89kd6GfgZddJ3+mNrPHsEQbHurLcRoiMI0vBRouqu/3xkA5TS
8SBp0/HVmK3L7PEW/KB+ZFuOMBLMdt+wnZe8kk2cm8uZTNPjfZEBp1/bXalh8Ew9lPKrLiSAk3we
Iasqs/GYFMAelGpirZj+ln8r800dTRbw79SXEdLRv9VeKv0CVHpWr4VvIalg5oAop1rc6GBPbH+X
xybVaocda6HcL5ppwuvKoKPJmTTxU19J/KRQi58TkQ8CQKWqoJn6BiDdvGanRdhWL53SwE+LXNp1
XSdi35GDKVlpCz7bKaEF+SmfGg8IEtlI/LuuHx+15LSwpidiYr1D5KmShiy+ChtrC3exSJcNaI7b
tBAUi5C1ktpRYEqZX6NtkyhcuhvN9miOo1NaaFmqKNqELfbf203iuzEmAVa53TbQOtfX+KSwpmAt
Gg5n60l7tCSSypXYeGM1zbxJ3S481hoCUppPRBu6RoyikCh8bt9D2N2STp1ZRB4pw5dVPz+K+4Cv
R/nRjz5JQOPBWeTP9JI0Ccihz6beusKGYxYyqPhhtqHy+oc5KGNGulAh3aSrx1C8/XYqBQGwQyiD
Ks1VQ56p/8hDmvW6euQ9lD7PK3gRkCYaVcXKCmOgRQcLkjqYEgaw4JtgS/SM2XIIrEq838kfmMGj
D4BBPIJ4V5TVy+DHukmj36jo
`protect end_protected
