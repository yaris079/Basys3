`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p2VyGK0MidyEAkbJufUZZIAApGoFxDuEKUDOXiPPP66aPwXHv3JGkBVyI5PwNK8H02vLsm2SqWfI
D/2YjfHo8w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YJwmwxsNIgxUVzVBJRytHdAscXgKB6Ygn+CPJM4C/86xOHDaCu8rM7uDddcUsrF2SP3dWVPrNfe4
LkL3cR2uIRItKODeXnuy/WXgPRkp2U3DiuPfbkMiEQsaI+4kZT0jgWi0C9YHxNM99yCFJqZYNSpv
TQZTr2kLkJpHFeD8GLw=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
km5q2kiKH0tfuOYiZ5rN+eNUkLNu3PZfVRkXPe+gfoxtH9xOp59uib4lqlMzKyfUwevYGVe+jViG
07ViNvkj7bC1yAZZbnENb0DWg3S0x7QnHBZiacjw/gSqrN6cudkwYfXqRThZnokDj1Lpuqu8ejEw
aBq3hnV6ibjeKVkkwVgGYmpO5cyflA7ZG82fqxyKBT9WQlOJqscYeUAU7m7vDqWV4R/iWAOPkSBq
srWYufHx76mzGzbtYOUHVcj3J2q/tkRRwPiC7OaLFvNP3aXiwgveLn+rGYWxHxIVM3Wqf61IQlf2
iE+6EVLzkKohamHIbV+pErFfnV2AtdfNw9yUPQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rBJ8pJaa13H+fXdLKl/jZy8aKlg3j9AVbJy9zheQN1C4DmcJwkP9nenPmT+jE4GPPVacV6p97RRa
B4k74b9uJ0DJCs86P3jBU5mWaW+ow5WM2uMoYBOwvRuk1bG+Nk3xsVVjPwm9ha60DzTEphCa0IDO
Xg8dMRE1iDV7dwrIw80=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AH7r60rsQSrnZUW4OpeErpYnE6vC4yjWOgtdmWXeHmiHJYo7kbDgyJ6Jun5M8fd3DjOr8V/TDdMF
veiUoL39qrBaM09tbB6t8zHg5NXzSAzjh7GnCmzB2At7FXB2vEOnXGr7TrGv+X+OGnX/FIDY3IK3
iL1YmQ1yemPftfHj7xeV/VALMac2prz8/P+VTHlsEvu3Ds4vL49RBl08CZBVqy5YRPazq5r+Zwcc
cgbonLPtNtAIuCoVk13S5fnfzQrn4fE3bjo91SnYlOM/nlmCh8pna+xg3jLyuTGF6wgIiIa1phOH
nN+js6VHDQhOBrX/iHe9NpwICbXSdiP1A6YUxA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 25280)
`protect data_block
1aQRvcjLf5aiBi3mMYvVefUBd8LlbI2stA5zEnG4hu6/Vcbu/ldYiRhRj1SbUd+SZ06Gx8Wx5krD
s0Ki0yCU3/ri5znLBB7f7s6/cOiO2V/dhYZUDeTCcTketHXVxfQ4OUfO8+oBGUz4ihuOcgeZhGmD
Nt4f4ja/ey6Ilmdsj/FzccMtu8rCTD8uds2xpRz449jNvLbDfCjp32M/pYT7P1hfmGBxV00+TSY6
YohKjihIXbvU02l7Ira6MEqFrLMTFd8Aq4Iy5deEGfadZTDXM2eDz1r1/VQEUkVSAj9siriEvI88
jYPYP2UGHKYEoushD2gGdQjf3E+bH6QrvdmGMg2ISZG6eq8VgjQHk0rA8NmskaVtIA2U8hsrsrJI
G9Ay6Z41/wGHMzF8jZaiCNbqty+5HNaaoUkDuLowgWYj6wGNpNw8uQSregvgSn6idgECDsW1B+50
jSwRzbUhqNyO0CBG8HYg0okuBYMZJlmSz3vJrVEDFmJTUffmx82qf9ntbNOFmKuUnqJ9IWctrFex
UjO+JMOzscTYhbBQMWJRiniaFDa6XYrnr9cJ9bcOOfHOGsJa5LKplJkKo34F94A8vt0H9ZHcY73N
E/MKsNQ1/VkAND4RyHGrZ9WGosxD5HTbRTjPOa/yalTD7YUuNEBI0Sew6EbbnmzXwARlYI4d4HXQ
DZpkDWVmT7DbVRHFii04C4zefiK5JlnIDe741oMOr932U71h38yjVYI89Xe8h5KOp2sdzkTjjQg7
43Y+18MK/kGeS+kzcCD/9Q1yXCnua8q2dhSZPHtVUgUZMv2A2wTwSaaYa5hrN/sBvQxybwNxfcmS
xtGO8ERwMGvvR6QSchfQteKLGa9r/6OOXtX8fztK2zYs5ImkmqQngMtzWJkwWes0IY1LDGfxfR7G
JD/3u2mc7kTeEL+Jom3cG1wRc2r1WkU8mJdG4qdJu/X99LiM7s90s/BjANKdUzaa0UsglQM/a6E9
6kIQwCoH+RhPVwJDOUmCh04eypm2GAf5wPYYVL35kVdi2HZqicAeuYJV9F5UYIr5czEfgr+KBA69
QMgsiZPM1UC5EnMm6TbLb1wH3mjBxBZHYKOAjoIi+EuF/YhoMz27loshjuzjOnhe0wmYJLkCFFx2
pcijo5CA78j51WoKO8acFo8hTduCCiRyGeoiu2AGi2ozdQL8sFENTVXSAB3HNGfxPLF/sMz0G8tV
vaGgGFCka1SuicIZlk5Ct+ZdfLCUaL7QnbmRjs91AFJgwDqGQmi0R3ZHEym4En2xuh6VhXE1XJXn
XU5yz1yXwOu6XRiUNZppFjB/uC/wU0+tXZxf7ztaqz9RZjmD1Wlm1wxQ9dN+RNqdHTN7KXJfbItN
K5YiuftUjdHGmKoP01+HYP0chr8H/R+M1MwBEGVqKLb7bz+w2Tb2GbwoKaDR5T03VW4BQyF/nm7t
vEJMFanuLy2gQnT5H6WXMAVii4qTBeBGEhmDsvoXhtrNB7LYIQbpNnlfBO2BDudtM281bpnpsJeH
MBm1dOq162V95a/cRfiKYb6AmBsyc9/9i0PzQd7/RdgywmBGBYuSjE03ajqdz4lsISnwVRX7kmkE
BfUw1bhIJAz5K6/yQvrxOjf7MRk2r1pZTMIO0m4gBxyzkANEJhCPCByd3tAsD9GAc9Ytwvk5Lg9J
tIzlJ1Vljrq6uEEqR3AK0YA1CSSmdhmnsjZcy8qggU1EXacDlJx3SBnnvG10VguipiLMXFYKZkJw
Gjb5kuVglHduunaxvtCR59AfDVioxlxqVro6R5SbuF7L94v9xhDmMcEH/DP6bkXUSvYuwTgARWn2
ssdW4nlFZBrBf66xczyXnB5k91cMNNcqgTJ0dGLBBndd2O1sv9tePuBZDlirS3HI3pYD0o4WVGm7
USAUohEyMF3u2Sw4id4EgyfWW/TzFUK56wkO9FA5HjXCU+gQGTI7m7gI3a6Ym38w6TXnJ3bLOxVq
YACL7uQLaFqHMIqhwNDMXP+CWk+Pe3KVwbBhROP95nlZxKB2qi97jRG3crZBZiTFTaqt7y1M56Ei
1tt8LECUmkRv6c028AG1PbEbQpX9mW10mq555iHbfJGZCtGG547CVuYE2uJOa/FnOhO47sVN/tId
Tm+fXJBXhtu7Xz7K8fA1NbZJOI2qDkclzOGXHd67sLN98K894W/y16H9YIBZStjahqHIuVgrDkyF
LoXMv/kkaRMmGDpKv/V6kcUEDTFHvBLf2DZpsUghk93uhqXYfe/7nlG3UhMrLz9OLUS/LYfpWEI+
rr4MU0Coeui/YwkLE3ncCatmm3oOxSF2d01JMNltfYS4qfdPy8lzSU/IwBpMlcQ827+McEgiKiF2
0dJrgs3RUE757ydEX8QaikKxL6XvBFHHANphM+E9ZKTE4Wylts6HtRbmHd9mO4h0sCIybXgTwe0L
x1OUUv7uPjq50rLc8DrhlGPBWWIx/woRGUGRGSEi7LxrR1E7TeN16x5Biv1zmkbHUoSXpZ4EU6qJ
JU68ZqxxlHR5RWLBFCuXdMkdtzSEicrzo+vgBys+e4ITotwvGZvdYeA8INCQMNl+YOJfwEUHaSAv
x9rfK1bW78r6HHg9HZMf2Za243DxbZPsn2EIN4TVHTspVHO4polqiXaM5UVfDa6XbqAHpREjd+Pe
lFeDPPWfthiVBsNmRfNuG0yTtPjCqUoGDrkfl3jnvROuZyHqQtCg1J1j3XtE8S68VSO5DF+LIQW6
kJaycxT3K5udiADFQJ/rDptDtMh1q3Lkd8Pv9Rbj9DvLz/+NXwAKAnWLI8/xMPIdtZuRInAD25mD
M/zszAyhePj/3Zh2OuxAeLIPgl4FKiU0ZRx8LhdVt7RkEXD8rRTqOaZtv/KIqK7eBK7Eb2tNlQL1
do93izFE7ABTesoRo77JWhI7ru5BBlrGVittXFwHEkWKT7fOAWQSKPbqQBlqmxEJO0zv/jVUa4+n
u3FLxBhyIdRtTgNVxz3byUAdfvuBGB9ynNQdF+ggmpSjYcF+AcXi5NvhznHBaveyGYdgT6LhHPyj
r884G6cfvv/rcOC+LrhWOA4B4aC/ydM5z6hEXJljGszi+QOy9cgOdnX2uCWGEgcg1++6xqQkK+QM
U5TihrZl7H5vbod3x0wFLf6C+hrD4iyrrmJgL3FWgByr2nnqJHFAkLi90lhUyBGZTiqJcEOaV8M6
RY17DVyMn09iDNy3cdZ5TKwBIq7BnmXLCi2E/XFJjykWOkYkVSElhJXgCnz00V3QqyA6siYTRT2M
/wlkWfMCpqD4LYAeoRuPrHoq6Ax36Au1u4TTLs9sy/QxacImTodUAlAgvTH9/c8AyIM8+oqJuMoL
DfhNaEiwI61ypjSiGZvlJjp+rDLv4ML1zxnXdNf/siikTFVDWjaLE8LaaAHPOfL20igQIkVxUxb0
PEHo7xpVFAaYQhG4REaO1gZF++Xz7OflSK3WstMc765tmE6nIvhi56Gz9SMLYMgwn/rtB5eRtXbF
Qc9ts20ar2RrQ0XzXPjn+W8TY8okRqRmPoh3znZF/nDsMBxP9HkqtQFKOUlLOxcygbaJMtW8soS1
6tU9glybruxQ5W/17jDdaoNNQ3BmYpQw+l31kp++KFppXaUBzckBDHkJac29BUbplx/ETru9F9IU
SmitxzsQPUJhprvV4b5OHYRgO0bmszhrJiKeRhPv+vpCJH0Jx3Ht5VQoZrt5UrSI7JMaKH4y6UF9
e7V1kT56uWTNBd+QtGZcI17av5rMYmFzcjDTcpjPLJ5GufoPvPs9sYWiN9ADqKI+daRkQmO5kQtv
NMNjcGPrsQhzdthz+uYVY52KJZGEsN9gwT4/igajkMQd+x2UwQ45w0SextHZu0wg3tOzax++EtDd
TKCo2hMwmLpvuRbdQ8o5HURbUJsbY8fklxHVrspu5W59nf9nfjZmRf035DFu870WJjB94ZFpGFZN
hPnL/HZeAcwQXi+U7SZo4V3MajTzCvcvhShZpOqqxdQS60reMh7CviaVk0DLyNv1L/EpyElYbTEn
Z+WbYFHAZGGMqKnaZG+1ivls9jImBZ4F4Y0TsmUL6zTCXA7V6GdaBjux2TkpBLshjGBfNhyYsLBD
tlIQwfSjACaKj51KyMM2PlXZ30hL4PLg+HammStqzenqong3zSBGNXSmdHtgbbFOHIjOgxRrYbOT
YvhQST2B0EIRynF8R2aVGTZ7WAKcujNJoXVnndlkIexV1e6EtBrfpJHxt0n6HEU+atsaBTSxkPuw
Fcc7pqenJ0QhVInA9M4IyrTFh3DjhmcmD0Q4b2t/d6lEJt9zBEM59T/0Wft43o9IMygxJT0Aodkn
feHDGsngtVDucPBWheaY6U8uImcRafJ1xnrW4v8u5CX78gPrgUHZmF0NvrfE99+1EoMD6SNeNzCl
FAkPRE/mhp9J5xDurJBxFPbc6CkfzBPlQvNQ1AMLOlMzOKprzuTOqO0F8QbDo8bngIwoY3dyJe4p
haBkpenlKm7LypGIipEiejvDkNBl5DrO/LJkoK4TUy0y2y05qm9ZFcIigSRiSV5FTQ1ADIWA2ovM
K7gjbsGruo9QBKny5mvfZ5Gf/wH/i1R3R4EtXKLjj7jhZbdfFhQd6nRFkJO4SeZlvi1u/nDg8Plt
6P5MZmjFaF88rAnCyPCruaIuQ4Dkt5m2wPa56VlIalbBy510wvZxrIfryMpE5+aIA60HZvxEAOyo
HX9NTUXBY686qmMimQ7NVWq4B6jiVdxlQObrj+C07Mam05E2C0Pb9vmXDe4UjGw/Gqgkcc9OCW0z
HJL2zOwESY+xIhM3yE5nlHS2pAVWydHU/5gHZ68sHEZcmGej36O5AYh9mAoUz3fCjE7z3Jquh2Ne
+L0HPcqFB1F18NvGMwczbLVgWb3doSYBcLiSvf4OXgzyhwycnhe0tKZtaI0fX0LJCVc96q+4KoTP
bQJWz8gIlW4tlU7QwxtPZ7j3GnlQS3oerP/bQmkcCErlovQwKWw/tCyiyCiDS6zeXoLYzgZANxlt
SxH3aUcouHr/HrNpcF9ggmepiS73WcxxTwatGHvGfX6HMVsByEDXb0SQAkak1cSZubr+rkNk3HoR
Z6jpx+ZHOw2CETQegN6iN3G8IAEz237KreCIg8jtGe0ytxb/kbtBN8dFI9nbmyADTI47EuTmAVg2
+jwNQBE5PAWLXXRuqWW13O19JZsMLVx5GrCrqLgqNgUOPh9tUzLzfa/DGuEUIjvY88uNzFjBTF8g
zf/rS9JANb6JWUlEg8ZF+Yp/qRCRrlLA9qGnrM/7l+gxzeUUgXPplw+Az5ONqpCExrm/VFn7EYQm
bKC/g0rj+9zk47fM+gY8pD0F3FNHUs+bG7e4gF+0xI0Z/rkLatvBpvvnLOQXsufJsJc30qubEq/R
Lu+j4SMvrh+J/dmKFFT59r8wL3IIFHKUofdQ4VjvA1etR1QRL7LMuafyn539tCFoNc7yAohz5D/r
AsdlJwkosyZ/dWICSc51OFqpR2RT4PnwEQgcHusLDa0QLmjVFTwfmi55L94dAbbHFF18wWiBa2jH
XpLAdo7tjOYZn4d5RmSCY2hpTODq79La8TytIA7c9QbqNjwI7Mh2LKaIwBQ7dTjb1hJWqxAIcugG
P3FS88aO7pl3yod3BZu1zGx0e8rt4VR4MLvWrzTLNN8neYdbcm3V93bn9e1w7+diZDGwyuhCgGBp
woZSrAk2SuzS60fnNDEQ01odpwUeGcJzGu07d5VdmRH5oepRecADvUR8MZJFO1D2MWyeO/b9246z
mVXct+aum7+IoYsbySpU0kmWyg89EPIcIUhDeAygHmYiyLUqa/+mu1MUG5IbsXymLoEXsYeTiGOY
/diDFbqHfuhXKZRJ2jeOloh25uDNK9VQqmJhya2Eqpk3eaXRPO1hHCeFuqyVQKHFwV7+0Yh7Ciw2
/XtSu68xeBgosuP9VRbneo4uGZThkXYeHrivYr8lCJ6h5qEOX/j27CDp+RzK1AMb/3jdOMoAK7Ug
dUgv+I//iGeu1syusiUGrwKQRQO4YhKh3in4ONPc2AhZDEfWACZHu3PKPQ+GoewEAqLrYG7kgPGb
LqEo3OS/Y3o3KOpiz7kTGzUCm+Z3yqGePgHMk0M/MyvaLjZLvYvchRto26cWK4K/9UKv+E2vyNMK
PU0l20SpcWpuf8KcWH8Oh93Mkxfo6oRdeoMvJTP82DEblweB3Mc730BYqo3N6NDLZhr7pAn19X80
oFyiJULRZl6UPgOajjDdGAemJEVD7jwm72q547TawPdjqA1cCeIyAdfoWpMQ2C80B+Ql5OHNSdJ2
d8WvCai4TH6FsyolkwTmcdlgjPTdb5CMs/tPlYjKxhE9YxMyokVkoEpGhXz99RExHVgYpOSTWQfS
hH44ATohUp0J2p0fsYSQZheUtnaYQPxV5MXvuorAFlJi66IVEqaqtZMT7kVO/LcyOek5ydo0HKRB
QMSJP0LRcRK9bdB7uovUVTzaErUBO1vEn/1I/JXXs5VJow6FQKDs1odjA4D7vg6ymomQTVipK0iv
rxYqd0Qh2wKPOe74fCWuYXd2POrmNg7Bz3/BfcG6e4aQTECELKhHko5+fECBEnUiPsdEmSaivXkD
G2Lkn7khWunXSBes7JF50A2r7Y4P73lDE9vAgrHuTacVfw1mztUl8H0e5p/lNX9v7fC4V+TxNkdl
uhasu8dIIVPijYQHqk5ElmaJosJtYMWjg0EuqYgdEbCjLEk/HFS8lQdnufFFN2o1Xx+VngJFZ0j1
EwYEQBePkqQgbAx9TAi5OATIguMP7w8pTlRYK1AffpkYOYKmME1TNJkyS/7tlNI56dOS3BtEWSAt
Iqw2ZOyKbRhUjNAwMqWnWQ6po5bfywPYgG0QiJrh8wxPFDVAS+/0869/Xi4llu48BwmMFs5Qr1mA
PCLaC9X/yQZYtMajF2uVfq9YCICHzmowmaeDcnjW1hJaWErfhWVrGgDSF1bT6xUQWaJI01MjfXik
SkLysa1Y1ynkocE6CTAkItG0SrLoaWjO+3eE/KxG7fpcu0U5dj3+beEqC+GoR4UaridYkHEaOjpJ
LBXv9VoLVsFUl4YeXcTWTJFvmmOuP8iEguToCoRkm347zMJ1efTosU+bQQOGX8WXlLbrQdDwBwW9
gmlMNK06wGzxFxMS3xMk9D/3Ojw4MEexApLDH7KatW4JyV1mXdRylpNvlfVt/R6qaiyFK81ZTAxk
0HQ5SkEpu59L0+OHL8qTwWJ4OyvjlgIEMTyfWKixi3N0G4YoQeBxzrvaLR2X5Hh3rE4+O/7ZjG1v
wTzMGw8BF3HT4yM6GMQ1Oo9mlNHbDppV1Fw4RtPIThmdXHanl6dTGzfIQ2iMiUMfxbLmeACXniCm
o+DGcem+1C3WoYY1hI6YBTkrY2i2jsbI5o9n2681P8nrDZnd09H91vqc0iybtJROgjn4Hb8Mkdvc
m7xwwpyQ7stPs7U8ju1OReqdssEYkWIYhy1Q+6VGTCO5R+egqF3XcH2t9WFLp2g4vRLaI/eeUULg
zbMBEvImt7AmTGVSz6PHa7ks9+KVfVbQA+WMeF24GMBRniMV0BREjwElFUqTzDfYnk7VB5UDySZg
qZxvItRGeUHXXOu4k5DLHY7cT2IMSL4+8rxYfXbRhM+rrEBqNJbGQQ+UB4YnrLDl+hXLu4uaHt+k
y8isZ7cOHBSNqTt4iSolPT+NqXxTVEAoE8/gpZ5SQyTjIhjKbvJC6jAG0iO6ib4T5CHgSpEitWdH
NR+oMDYo6O+btxg6U1OYkOD1EqEiVmBWcWZU2KfzpibLsULaI+c+gVu7jIp5NqkcvVw0ZAzn0i8P
mbomVJBBZzGaFCM7quPPxllykPe9vXOATfz4C1HSibfd9/0KRBXZ/y4jM1g+PGeNsT38rgsdfSV3
pFMrkOGlRKwyFXgVuFlxn1LrW1XcCXPVZRKuR4oo628tilMxJA7n+8WDRFagyn7a7PJHaEX3fhGe
mI5F2kRjtIozkTG+h/e3Wa0z1feMf30iGwZyFq9IIY3iqVH9hlnCnsmOdlsX6LtMVp8u8atis0S6
DPk0mjVKCoj9AL9e4+lP4E1dSa++N1gU+u1CAYJw/gQxlxHpCSNSc/HbNy+WyAbDUSiQN1Z45q/c
Y+idCQqUBgQVNYaPArteoAs+HHGTubF5fpzDJ3Z7SZ8317sJXiAEjOeAjsHQabffoj2BsjueAiae
PeQAwa6I9BSwqvXX1JWM9wlc9rM/IWwzC32x0DhFQqteqAXnQfW4mHKAlYuBX92/e+veOIXssVUD
acPqiYUkmdW6vKCohELR7pUOJtc6Or9SFVtAKRHpsJqMpiqfoV4nFHUAP+o7czWFJawIAm2A2354
HSyQraY4aRBEPW8zHZjmefNFpR64d34yCFaZgAf1GXoX9KNkHqa76tD6wb76hKSkHx2bSIOCK59c
lTC7FYjlRsArUC031eW8vKEPAQnI8TUUZN5IkTLbvWi4U+GVN9BjyoSISO1LtkZFSgOLsVA5FNVc
bviJYz5aSujoGuI5nEX2H4es9MK2oGwbJEcx13SDSOA+9NBW2ETwk5CiebYTq8dgTRB4HPiRtHic
N1clrv5R8IKVudX0WrobqdKiyPW4sLQTYwc74bYIpbMgeHdkWglE9u5ieMf64Bgwiie9/dz9QXO5
NlRLhlJSrxKiFqvpKj6kzD/Zb50WuFsSthin0d4s5oxnPIba9IPTz15CfaGxauxjxxDaQgU8jgot
lZM4gJRdWYZQno4AGW8UjkvJF+eqgrGTMMnFnnCcXEUSN6bffRzUdkApB+tvKiu9zsIWpTfBbgXi
mpQY7bKDy+PVlOjVVmC3m3DJRCNtsFtDE6kk0p2a0xg0/L1LEeojEb7/feFoT05N7g/KFY/+5yuu
VbWpV9ORwDajVQ+3BUSxVD91ebVwBd1SMe2++BQ5d8Wyc0MFEJJPyKzedY+QK83dcWdGlIzwenoY
sIHwr//+4yx4oRp1XSSSpBVzoFFZ9tLG15EGpUdQqjRu3Wdp4OQeV+jMX/D0zIEmpN3mOiWizSgt
5Y//Ktetmg1c5S8lA+WVLVr39U0DHGbW9+c9QU/Y985EVx3k/NQIbXGHdh5ahi1NLJAKozaqO8Wf
2QpZ2EHrJDsUMzVF8S13kJk6CBj4OI7sZLV/4lQCbAU5zzW0V8skMx4xGm+fO+R+IPq/z8b2PMJo
bUP09NmxlXEpgXSwze7DIsbohb6efxAOJNi48fFAb5XfUDBf/wGl6hG3Wq73VXjDrjH28oqwlaQS
5EVqSo6+96h8x/c3LwJPZZTR/MatmDo1bSCnh3PGRzyTdHmg91BowTS2T2o7+glxlNn6SyT0iLCX
D5G9MAi4bWT8pK0foDymtp5OcEenzjJNBe5PRfmZIg3jtUN+a7DaOX7Hka7fYh2KIyFWJOXrzftC
FxzkxtsthcKwbYuOr4H1GrSHachsjuWeAcQ/sYytn7ngQcy5hiEgPk9k/O0XHzzUQX8XsVnFRjSY
3vr2FrQ6kvL4iZr0uOXlAPj003qco8g/w1Wmfsn4pFvq05cdPvyGhRI0Qk11Fvk70Vv4iEoe+V1E
j6GdAanEFvre1zSN0A7Vc4JTGGZfYQY3+aEmcfqwtxW8VObFRlvCK2WAvBVRzjfwoFguwWxreyLa
WQGoq7gcZUG66jNspN3RnuYwPVmu1KsPHLeyTx2FvbXQR0sF6Jpu86Hr3p/gS2u70Ot510OgPCSw
b44RuuHzjANu2eqIWLF8/QWtQpCbd8pwRrMz5KSBqYrrUYHfCcC2c10kpI9tE1XcdNV1qGZ3gf/h
LMPogd3iRuVtgZuDLWI0pC1/97xBVI3klZxorZ47cLMbplyv7XLEJZgsgDl2V+meLVLTTKfz0CMd
pKW8NdqsiLOGBpUWZ63NxSiQ6LW450ftrYHUwwiJX1Wl5wv6djVnS2lWOn0N//+a7ewBX6NfrHW0
fN5rL4MDwKQWRBYAvlP/Bj9eKJL6LHXaPei+T00vJGUkFu9PhemB9ULvkLXey0/ZTI1RNRkKqaKF
mEOvJMuTAxYdZbYq21CVHoCeCh54+d+/p8AinUqUQ+Vp7JXVJz37OQjLHWaxGuZiiSYGzgDuN2Mu
/HRR3AmuaC8n+RuTjmSzQylLvjfDNsfC6syTLlLejaRQN10Hprii7ZuJ6V12AJcnZB3dwdxJCNdU
7aJiz6zo7+HEfdMKNASUowmTOPnZ2VVLIp9PyV6X7IkFn/8+JYQnn3A1oxa7XeAV/zOFfTZsHJUw
RNPtcJA93a7jlc/JxVQK0A9SSMvy9DMWto/N44enaOvlTLAoNI11jGab7wkeA/+N2mfRGl/iIjwI
T/DdEwCmoQTrOsst2NECY3UsG2D0A+nbzGrBMmSiA1VrvkKFSxISGeD4tNKJB6SqroH8vgKseu4B
nQzwjFRtRtY3ibFTJS3Q5SoI42n7GHHGVWxBxOguNzJdccJIaNRsgnamuI8HpWELcwzfCYmIYz+n
MAmVdSC/JQS1a66FYg7MElZik0K2VwYmhLQKQ4D5YtZdh4HlZJOBsKH0YYZjZGXug9f5r72MhoGU
YBEC6YvGu9MmfSNXR6QrMV5Y1fSebks2/wjFq+bkLzCl8RVEtjGDshF79RozOs9XEYZ1RK6yjNq7
TINwsHkMWjbkEbJeYrlxK1sfk9LsKiYb2sCGOHl9v9FZ7OxL0HK+EiyPSwi5tFXZ6ZNeQdRE6KTc
pnWSRLuucxP/cmgvkiMA2TkuD1AXh3VO+t4CAexT0v6Xi3zbuW6iwdVMcy/LDlTiLKTRhuv+JTU0
qKcIJ8l6cwtAklwFsjUXp1co7cNDi0pDN1Aq7jvLukz+UrOW6TXosyGLVhAhrIgX/llT4gDbL2rU
tgzYaCL81w1lJSe0xDKdQiLJn0eM8GMVPJ3Bx0z3/18Fh0DG7iLV/pMJKTlluqMzZa/msOl6S1PL
n5MjRcZhbvo7HrskD+rqTsAIxoxO3V1T7h53x3u/fIwquDajhUbavkPRoZWSUClbllfTnEaUrQuj
1+PXfcSFC6rz3kxd3WkUQ25A9i3QISt3JtrWe97WWB2ditZ80KpozEP683xi9oh22HaW/8WDGnEY
f5I4TRiIlS787e4qVAWwOFj7evoZyrER2JQYdxnAZSopNAdx62qudjGPtAsShlJZL+HzB7TQqbKr
PkGvcTD4EdJMLoSKAuJOk7zXSUP+/QNd2aBu+qwN/yFTAG12vM5y20A30mROoFwhlg4m2k9HYm40
VeKjulDPy1DkHtVo4GJYwyFDRuajvBTQzSNF8Kfw2vSFDzNDy31LcgpZ6lDTqLmel8m7V3xqTtFn
scO9keMFUn7vwkSkEr3nHQMGmd4W6OlqzutdHgU497/zEFkRniaRAGnTt2UoZlDIbsiptH3uoBrq
r3Cu/+2IrrlbKxgE/MTJYNLb40KPvBOAdvxSFhQ5Bp06Rx5oa/PDuXvSu86jsNuh/AwsJi3mS4qK
PBz/vnUCvLx7IScaw/0z2pBKtFsLOeqBkKknuNiyc667NNXwJYAa8gInT+M70gh4lpa4xu187yH5
//I7SZA3l/GSmoL96R5zhCgBJgibGUx17Q0otXN1GtuWH9ZtTNrDKlcSKc4MglmU+og5FxuM6Z6w
Uh8FgkK+pukU7SD7R7TRiAvAEVTSdtO6l1cBQ4AZSkCADUDqwO6LHattr8G1l2TA55OyQnk42ofo
At++Q+t5Lxy/hrJiuQulSs6Po/ZM27RWmYX9+PCMpb4a/9C3ynZpn9l7ip43YpxKOCzYcO+jkkVk
m6kAAX+frqNaeJyEdn11NKsryckRi+85ilWQdHgcSHOdDL5rrJ+PonmkXkNC+PcJQ8cH8h1NteAu
lj5644S9SHNRAmW1Ajmy1Ym6gLIuK4doT12BkM3IKc/itL+Pyo6JLywfWYOKTkxd4bFk3wdrvp33
xGhM0Rn17oq7+QJGldmXm2jmJzV9jn/2z25oqAR7L18tbVfkqtj5UBzHPofh1fFnIvVnnx5iobtq
y3o5nLsuU1meiOh392/9HYwoHpPKwqo2MwPpxXbs8RXtxQqcXKZvd4bxdxf5iv31wsbhhl55odc5
9iiz/MR0vv2RuDIBTObgY8chwwNoRZxfqII3rJgL7xZg7njv/8aiqXo1cjXwPqT56YT6U/NZ8Isg
Ph+ueB3DXHsyuafZopNt3N5MrXVbL1UYeLxohatRVggsDEdahVqGnDnF8/ruS/66LOkc54RhSV6C
6I7HXzHYRLt//9JSwqKIyz4jW0xWEdK0zJoYMubPQ8nR4MiDBTQuG7vdoHUMzxEo0Xh0+tV405yB
A5UdyJ6e0s98GEJhApyqDUgSZhxv7NMZS2BAj7mKQtMfnO92nladcwTFSFi7/VCqhZFFW8CHHLL8
lhJUFKskE/Di6JoPil9OICCRyYOVuAztUr26kkGYvPD8w9fCvRDl3FEbF9QNrSTXpshtF4EVnBfP
PDGWzyeeIrHBxmblMwG5nodQIxwnrL1sQhoto1U/vEJvogxhWvDk2ock9tfx6DnNJ3whum7/6Nsb
L+VDLv9rF85byyXnHq3FZj+ZuTMfAKlYluScks5RdcVqOIXcEfne4jkYK05iha8yd/4QME2oHaMs
RDcqrCZT1D0nTRUCVT13pYvNQmd6t1A/i7701GCq6urVQ8MZOCyZQYLqltTY9A5ZCG5+MWwFfhiV
a3xuzTGnUbG4ALQQMUSKwbWKr73YLEO6e001N4IuMHM9ZX4aeODMBKl5hxjJ6UqTC4fogFIeL3qg
3YAd91xnfN3NxByqw/raIca1Oo++R/GzMDfDxSvXfdhxCgfURzBNAGWHCS5Y0bPsKpripqXaKS3+
RVAEIivv64BwOkqB7MAt/tWQSMxylecnmDMHq0T5jaPxCGwMWZuZ6AaUukdfYUklA8hvLrzRbp7O
PJPSiJTG3zFdLLk6Ujfmrjl4pc2d3sZ1wvko+FImMQdTwnT9SkFbxuhkADxFLugUMygvvtM8dAmT
Le9IzY1MAtt7MRaeonwhh6GoQvBydZ2sST3KVppF9GA3FXr3iQIvSWFWnKsepzDMDlaCI6kyc5vH
5XHCRcNPFcj1k4LLOYN2qs/2SmIrO9Lx2h1zncb59ZH7gCBNC2AMBHrdHIUO2QM70sCeW5n6N0ms
O4X5PUFJfxTC8KXA1mibAWXZvMV5x42q7j4i8TXVwatE12fiVm5a6D1C4plR58xFgztoQmrazJJb
D/8BAGY6qDrmStYCOmj2SHMWIdDqKzYP1bnR1PIFcQkbmP+GYPsLHnzhnVGRag7GSHDjOqJhH/wP
Wupk2VmRJUZP2QjOyhxMV5PS23vIubPiiAo7lJ8ZIl/oQpr/KSl3Gc4D2T/btL6qfvvM1KSuvP1m
khJFuncbNj1Kd4vMvriyQf3MDYfbeY9eXoAMhStM3RS3aBChLYNxBy0zm/43T38ZC3IO1kBJiiAf
oQrpj5FknrmekH0Fg2no94ywEGlEWQkT7FNcjpGm5UyCx/frYWH6iysOdkmbRD3LGp31jZnJsdao
jhZZwNwaqjKCm2TzA5nolsRhK2j4hDPG8wE4PkcDmGpZntQMjlFYUuPA6J4W0vm8ijEiIlJ3yFdc
ObMVMgXb+81IuZDcFi9E8Rn492xhrOuS0FHYD+0/JsRE7+jXKXkVzPS9Jrc1Rl5R0FTNF02Z3s69
9+L8K3n48P0xjEjdFE49FJfXM7Fwkr63cXyRl1jQq5JNP6ZRHSFyuLTZ5CKW07kIyZjPcezPZGFA
Sn4hv4kv8L9bvHeidD9fzLa5b5xHFy3Jx7XBJ5V+BLlSMNj3/jClKLdjfRygSD6rZueJtlLl/Kr+
rE7B61ABN2Sm3rE8QLC3hZJIji+JzwRHZre1zQps48yIgSAQffSqpoFj0K461TkjHxz4CeYs705k
hCxnM2Ccs5yiueKhVDYcILyQIGDl+f636puYx18OmulOaEzRtUzxlp5L9+/J26+mMW0UvtV7QF4x
6cuEOK7/Pm4UVRi1MT12jmC/SRGQcsk5WtY3tsnGt3QEYW9Tl4c7ievjXFIQGZ/ZLEht3WK2hEOD
sJuxCk4AUoSPxjOIAb0Z/LH52jxvO7rGeCImQ/eD/n/CUWUNRi45uMf1EhGXhuDMsvolw7/Dk5e9
cXYmzeJHKErHXDNc5Zj3Yq+FE8TySMStfAXK5pKfXOMmFkKpVIg0qJyRiWp1Ki05iWPUVHeIoUjw
jmu2SEEg0o7OvH19ln67A3XWvLMa8EK22sb19EZUJk4UzDojr7bULlWDS7vDdBpp3pSIjDwMXaCT
wCG5vTa645v7ehE9KHYU/XdepOhqBVQAQlODf0HKQo/ipuz5xXmH5yxDLqS+jRNYGxN9ERCoUS0n
jS+GjFNdid2HkJYSiJrtb6X/oFzTsMZgK/u/fp3ug+8bmpEkN5o9DePCfR2nq5BFhFf15uLGk22m
11syyt5l7p2Pki9q9/neqg3jnkV2dt8Dl0sBf+3FCyur5VuQobspx/V8mvc80aBFPUpdlgQCtgIm
Ei98KLWXOtm1POqobhr5l5wS8+vytL38TcXGRKbiAX7o+OWLP9vikr/cxZd8MRPhEk+r1PVu+wR5
tdrMpptgUSnvBeuA3EAkp0viD+YBLOLwGc5iXEsW97AgVZK5Qj8uGGWEXaPYrXlC060qDeH/JPEf
WHtPpe7LTpA/qnMSHJWPSOhCLcLABcQlmGum2nVld9OiFJUengUXQjOvuJXeFZresKM7prJmNyH4
SzTeGQUR9QOEoZLHg+QUYWlc0JtRdl3cBZ+TFOZ+N/8Y9DcIGz76VxhkVPzjfrPPdrXvbAiosw3Y
FoiDTpi2dcXA+33l+X4uv0MF+UDbdSHX3SL+pg/Pg5rGJiqwN9RenX11cWvHDxCraDrT56oBPj8O
cP74AJLjREUvcb0YoviV3lXLOXvyziz6TK/uKhDGf+WIRW9+Q6rjw6qnq2X/ukdMZbFCeLXEWjXI
TttSNWbW4bsshG2J9S4aEcy/D8aIZZSG4zy/h+GVDFDbbhFneNcZJrOi0sEtQS/VkDf3YwTiHz5w
PQVhvo+Mp3U8/dygzuP0eAGrcaT3gdOosJhlcl9zccki63EniZi1ofKNInrU8osgfdRHT9BIaP43
ho48BwNq1Z2rWweOGD8ZiR35q38Q5ebwAxeQlCGVwO8pbcq/NkTWuPg8ypukMbYHiOtfxqeOb2XT
lzDOhwEb9qN7a60tHQo4d3MAiyPQUJmX8gq7NfR6zzQSvbiSwQjqM3OfvgFqyn2TKxtnCblKNWGX
GYehX0IEnuLBKk9RAiXmLnEz+KVAAfhqmZlctxQwdCLOw+TN/zO0r+QAhZRxt1iJlkp+aOAFciPw
REmC4RUmlouhnehaC9XrW9rUmnOC/PVtyt7Q1DWEaxU+RrWBPE7aauchyO8zg9uvfQkdyp3uMTV0
jo5gZ7v+Cl4y3J+cNUWtgwGnZaBVOCwAqIqiTAEcmIKqQUWNzRLHveGUNTaeLWrSMDaFGPXC3PO8
TUtfqmztBo7k5mVgHKToqGzDW84yOw/Z7WfgKLPRNvYkP7lYcLcMhD81RxsOe4JqrV8+XtVyw0Bo
iDsrMMiwayW5Tp/VpimnSvJX5Y6WhHeeQN6+ugK27c/BMsv9BT7CEo8FysBn/Ht5DjSvxa0WAo2V
+rRl5Y/FMsanR3+GrJwcJ8euCPreTmMyjHXf8lcmKDOdooiuC5CantEPqM3kMqDCU/p8fAFlQh22
8TGgEIxZuOcIwQ6OmubCI5ZabqFhoXq5e0kseR6ec59qMUYaDaK+O0ahnOn3KYRS1MB9P0hLTVB9
CFw4wSlzdGhZGSKuc3znSokUIlnhKupMwghzWKMEfLIpiOSuGOCA8n7kv9Bb0T+NkkqIQXIHQjGm
cHVyhRFdhzyvTN3By6LRMVciaNDqIO95X1ACLLoZPCgZO6xHoeJ48jLPaOHWSbKkZ6v6oRXL2g7z
t38bBwf8SMeeCp0JDnkrBYutQLWtl4tq5gdhzMf8tMziRN8Kft19QFeZ5ZbxOz+9BIq85hb06aue
L9xAzFOQF//3fe1Wd8uZSMIxEJqo2XFpmKPZmnMA1IG6nrjHrr59ggBwzQGXihE55Fpakq701FLM
rCIdhp470lchGkhaDVsvNJw30H5dbc41XJTkkGSThIO1GBsczbYyZm6Af5R30fos8HxXsNHtgOLV
w+1EXCTx1mRnoMKzPxJFGEp3MFQl/Iqn91GWxbLtGgAQtPbJqZMMCWHeMmImLJHa0q6fJ4JVdDj0
3ahe/Vi5gMeGbH/hrwtQmct6OYQoPsfT9s3HSDCJKg1N201yJoB3prIG/stSNUks+2bthvq5tlNk
VGNDvu4cFVJflAH4bsLf8Y1wSLIP0r3DZc3PzMrVaQPPO2d4NZ79OIePhW0oFS/Hn2jrLnxElsZg
Yb6Xyni5Oo5VzIcNKTCNT0oIZKLacjg5D/mX2MUZF7gY+LjHil1HEoWwbVm3VWNxEoS0NEZFeFTd
23t2LAVCt1wlp8PI/fTm2s6+/DyZuQMEkUidTSv9UtAaJ2LmcDr+FVyoS4L/W8Lyq2o6Z3O4+DyY
nGwkO5B+SGcVQ6fRKQ+rqqJr5LVAkbwst4t98ySYU89ZrtreWRXKd/eVC/fC4uCY3ys0p4P+6SPs
QaVVWdsb1oRDXy2+nssRChMrXiMqhmQqp3CS0So5mavHgeRuv7Q3UxKlLWT7lNVKaa8z+djNAJDu
n5BYPMmObgF+ytDCumcGIXUqdPZ+mXSghox/3FkJcylvzwtnR9KXDV9MrS7CBmZiFzfo3atNPHe6
ask04wdNr2m5+1L1GrNMO4IdCh5PqZTZP75h6M2G4aMTh8DeiaH6dDe8edzIxS88BriEEGzaNiQU
SqTEVDrW3OpuLoAzQM5/Cynq28StuZfg1ag74UmUbssHXrzxc2KsVxs3N+DP9sXDjhPA2p/BFEp+
dNaL3V3KrSrOK9H9BN63783t6Dff94TJtj1R3Y8am89ZkkeK4k/BVCL9hVvdrPXCKlZC1nJb/uZV
HR4drje1HrDcT/fuv+MsCkUMy4txsbzfW9RcQmHEaas6LNBgZnNzNrmnixeEFlNJzo3yA2NMQ/xB
8z53Du9olkn3hSeXPF7eoeLVrZieDjphc22nsPWqHecAVcSoRYitCnZ3aqUcXWrjTLxNO9b/kGdP
WVrzCZBm5dDvDgueWQm5hoPcFG3NoxDhyJfyncYMCEPniXxnEd/Q4P1uPZxZKvZbdwc1PShuw99H
crzjzy+l5o+nDiKtNzGkloMiRgEbOFa5pyChVL4eb+FzB1yFeWPF5RK4isq19J7/TfjGj241md8o
7iYLHv66p3QviMpewPOOrm4yKrPdZuWVMQXzldyDqqmSz5iXK1Ppz0u87JbMsvOV+PH7tVHkzCHA
l129CG+wmAhfW30LiletRgMk31B6pRVqdku2taaUydNlWxbYqdQ0AFury2GZwxA2IQLLHhLo3K2H
K3mu9bq060OnfZe5ktAliISw9DEHMMB8Y1XxTWLmPZMnwI4Y7EFhYF3i8aKuBTzI8OVpcxgBigLK
T85kzifAz6Z+MHp2S7AH3PkMJp79+V+7uJurTyte0dfGQsRXGuHLdNw3SgkaRG3Rywgj6YpE75vj
i+RV/qiyerunoCAhdm1+eYDEBASuv5ReBXLGPH1fxD6aIkaGfHwSrMudI0cf39P+Aq/xtm1fAhwg
MIsc1fjr0me1qsxgzWW0d4DpXh26oSN8pKYNWRlZVORDiR84ZVEkbQL+cwzXNPJNZe9klzF6aVtg
B2wrjDRJLDEYVChDQmAFmW3TlkIyjnkmubfIWw5KiZ5u67c2upGjC4JYHSov+uA4Iz5jM4lxMNk4
XmDasfpXuZFED1X8900NOc03SnYpBxaqBTx8T9/BHai/N2XlW2ev2NK2uyXDYgc6lvie0uuA7G9V
Zb0eeHqj0UfN/1ZHfoc6IgANhLMOQbDDOeeEa5Clew33gg6qC+mm7l1N6r2Ifd0/EtHyllajMlwG
U54M759aa9qKLUNxBtaezx9Z4i5qjk1tzYCVvR/ZTatvLiCdcrth2AdAjLApqeTNC7glq/aVaezQ
kSH0qxwRBFyzVDO+TCvoiBpFw+GE/80mV9PQG2s30t2fFJS/IqeZKsA0OgDp+jLaAnP+9OEbfmZO
Hjn3xjL7W3lMIuRsn/EPwk3C4/OvA5RU7v665aurCCJwU8JTvGi6MdJ6CcRequGtln2TgbZiqfmb
gYj3aY/Vlly4IB2tQHFmZ4FzYFSqx/9H3R53UrlYu1Gc/CJC/CoEKZrYDdFM4L5pD+dwUy6gXWRH
Xf9ghXCfVnpmfXw8EazeIbZt+EkPgcpTG4wBZAh4X0HHNDClkbMBACXtNNd6xUaMgAdIs7KOeI5G
+Qda/RaLg671sqdcxtLPBubgy+UhDWMH4T+TumtSGQ/NqI2rfNeM12IwLA8ztALI/tPTlUkQPQaG
/57r1RXsQ4MJ4I9yPxex18zTszyl5ieWu7OTt+QSc3RMd+T4YinCz/Zvzqg1EASTj3K2nN59MCtx
bZmepRJY4U1LmySNoM7itJhDBKmJ4yrh6BGwFqMDd15nqKGwgvUqMpSEg5hj664VIqm6hwgyA5+B
ZqNDfOcXBB14p98b/qo0XyNhilxwvun1jac6lmlCTNrSzmDL13nMpsWQ1Ne2DUai+HtloSRX3fcm
yXJ5ESBCGLs1xowLzO0RI4qZaKTHGLOkaHmR0RlBV/op6AGRCoJWjhl3eNhYFxQzkqvWcI1548ws
/+3byEQXblQwq5dU/I7k/UiGgEsN/URmxAiIu+oAC2PQhFC1O14zZasXnot0rJympHSDNJm5KnUv
OGahMHI/gV/7i394MMg3sNshO6xe5tMBrPi/zndoGrFwUFGyFhRfPHmkgI6QZ5MT9pdlVmdNJkni
2mB6gHegcwJP4+H5Yc2MGE19RBxtAkb1SctrIJ5iknkdbyQcBg0uTkuK1QWxxiejaeP4T/W9JEGl
WYoGE/meM+M/CCcSy8Fvi+iToEYHGgV5oqOV2LvDxaVIDzL0/Pp0VK9vP5Spn1+8UztpHhZ3nts6
QU4Ji2hksysnAxj3ZLK3nQ8ugYKYcuy6w42M9bl/ZfiVkVZ7nHs5A8cyDPtV6TFm4/0iUqpmtcoi
eWxjPa3Uo9iZbDnIEyxvRzsWY+KgWmc+dr9GVD8eDX02Y0kldrsDaGYhQsD1MSBTdf/Kln34lFzB
Lkcu1+ZirTvzRixrMC1u0eHuclA/5WVKEZ2J1lRrzLnNMB/ksfB8CqEduKeGvx9fyZZ36c7hUO6c
NUffqHFbn43h6i4Jmsqo55v0M1hq4LuyGrSWL182TR4oZe/T7w74dbwBXPeGfr7G+FWXCnG1W9l9
kzJx8XUykKabkU1fBJvP4L0W7JXNrCWwfrL0Y1pOOm3DCwJOwHZrJ0sQPCsqY1WHX06YXPiAbvMG
6fbEB2AQqESwMC9gDrXky1WmKLE+oaUXuNpTKqhU8eXYofZbPlCxfY+XmswUXzhJF3UWBEBNAgCj
LxrtrvIW0X7NQA29ZPENrcoR4J12MvDSZQkIBoholZUgofdKkkRby+I5hpDNp23yUD3ZQxCaZ/pK
JeQFMHKcZvOBBnAc8aDgbAVG5tzvgipFApYcBjic4E1Z1UkYc9RbjmRYa66dgiEQtsdkO236t4ru
qwM6AZ3sNaDySui2bJvYav7huFLaaf7oO/DOneuEIGbnimmIT0JPa+hrJaIxqFKRa7aKm0Gk6Kc+
8elabcHw93cuPP4N37rUn/Mt7VmNL4TEEGDHOgW7iW+gX9a8Tup/4CoubgrDEFXjdZSQMFNHP9oj
ETyQPfvveA8wsPNKXscvTHBAFW9kNvNDoU/W208SosIhZqUMP9T5UJLbad0DXZd8Y9EeZi+CacZ0
gRf6IrOLmulTaxPhhNiopXwC0cjDFKeaPjAQJ5HIQ84w0t5jEGSs9mirvEj7G6wNbQMcgJ9PwkN/
HjjQG0OMHW184ZJp44D6SnMBIXFu05JiTPx77TGtkTSYnAq5wfsE0dja1gVRK1oOavDJY77r+GYn
FHWSnjH9qtQ24C9QeCQsGn0b6bjhwOYDsVXnMwz89k48ZoV1qV6EqnLrf8y5BeSa5aiXaDqsQ9rC
L8y8JVZDo8Db2xXqAcgTWjdaI/8vVcLHiHrwTuko2cGxJjuxfEwwmYkoT0ZvKQ7cCFZQ3KGTkvBC
cb/ecIBQ8WPBelyYNQXJZVf7gdkEA1Qauw7OgBXzGFY+YLj8+npPd4Ay8wX+59PJsVrUwjTiIpB+
V8rRO8OGJe4SO4o1WQCUCRnS0UDUFd2sk8s/Egyn0yOvnOyTukWYJVYU4O/507gMDZbG2hqc8VBz
mw4b3qq5WTMhqeWbm0U3rr1ds/HfTl60SszNtmtuF46LRN9sMm8aLB0Yh5zb1wDYXuiyZdyWltn/
Lfg61h8WMHrAPZfw+62uGEe1FvXVzQ1ocJDBqsNYlNgK/bo9j/jfmSkDS+QQTkULFQapXdWyi59P
kkUesmZgJSV13gJHLCAN8ARy4ykrPhh9W1Hq6jWxsnl41SSrpSEzD0LxhxyfJ4oTzeW8TvxqijTq
frt4w10iO5qn+0bLEWDb1zOT9MyzHBSMyhEF0wU4VTIEAdmRRKOHlN3kSxBIucFI4Cao0vNYbYX3
fmdaaJ1BRrnZX6ry2kt4Vs67cTt2jur9CYbh/wHP0j9ElTZM9KgN6LEYpo3ZIIOkOU3rx7PYki0B
SvEzkSRSzhUEqt6QjVol4JN4U6bPYa3T8x/VlzNDeO2XQvC1Uq9x3GHqODUP2+TXCGLifKHcCCaw
jun0GXEns6MUthuM59TZfDAp3cQ5dnU/Nz51z9ZKxIojnEQDV0iEisy380eI1mZoH9214sDSnJB/
u/DHGsBNIka17a2MIwhswLIVnQ4Tx87ZrETL4WmuRzGhA8SvQuLbqkwcexThyYMQFti5GyJNougO
JNuqrRCRhz+q+ggc4Ela/mOIKK4i4BNkV/6j/w1uwewMVnaAVx42hMk+t9scCVQ8+WdEymMNdM2F
ifbfw97KX806jUotQ95vxLe+qSE9yAskBCgjp6XvdXNviw3lCvM+M+0dLTvlHKopVTGMvDcUdUky
U8gLhKT7brZmp/I6G8GMq1fyVQ0asz3vZu2LuMry4WrLLxwRRQI6aPIAhTGgwKWLT7g/uxXsCnqU
E9AXR6aw2oU0EqTTOLkNhij4Gg3foqO775dXvLpEcu6VhNtCVcXT/hSoWBBP/dFyMqShzg2Q6NKf
NTWpwWeBokaS5d6s14u2V5JhcU9sZcQWGdgfzxw+lt5ncycbXegIFeI4/o6VUUwTSq3la6ED0y7o
vMhZJ/gfywKT06kc5/5xHqNIZDC2b6TMyArd/a6GS2mnA/n/hs9riUCN/y7x9TeTDQjAW3qQTrPe
sqLWTrqnN0osM6YEMbLBUp+cZTSrL1qzGZfgK/dadsnQPSndCpn/oScZOxPzkGbVEM4lA0s5mClh
Ur9C+C4k8QMFWHeymkfe1YNRWrZBxm5bTaIVoaZEqjK2qxWMfaT+ZbDd77Ox0Afav/Kl9+vqj40P
s+2gXWOj7Rk+ywvJK+5vLuGJ5MEz3Oy+CkeYzRZ4YFbqZwGjGFSXF18p6nzA7dnWACQbh7C0o1c5
J2nEghQRQLUb6Te0ot7ZrYvk5Dts7kNsngv6C+BxWVyL8qEl3h1DKgctAtV0ab1uupVNlGMmTgdk
DMeZVzRv0odBlEem/AAy8ILE7MMy3Rs5vJ3Ys/2rnQtQeZxOwRl9oPz4mR2W4IB7uTKw+EOW6/Ct
ONg2UFaO9VPo8v1pQ7q9vzv+1rUgSlX8jacb2mhgSklb0EAL327Y1kHtZTrUfT/csFTprQO3oWKH
Z26jzSERD6Dr4XU/EN9zj9YdUIutCgwUmgFXx2yP9YsVR3UvB1mJijkYN2YUmtiTtCKMLjH5VQhp
oGzq5X0ZB3FJyYTrWszP93FwgJT36s8I3JyGsnWwA4Zo9gx/1myQjGmE9kAbHtNeiD+qgPnbEbyq
MK+DHv2Dm25cS8Fe9o4IXlB463cM0VSZ6Z/KVJF2wSfrvYJIWbnsCl5VY0yzLlwqWY2U3n7PFrw+
DxQehNDeFTKaY1ynrjTiyMNL+34q8d0V3mb6a+u8yaG1TfMiqFk7SbLJm0Le2/s8qfLJfTq6MTas
76WyP+VJRx8/CRmUiMYcGCJ02YTE/oEDKqAo2buukeacp2JBunQDnTLfqZMqCs9zSPZZCm+mzZhh
oQwVVax/E6dBysxaarLvYBjUr8DOgD1EdQCmFw9ZFInZyjC1asA4almlrtlhR3C4qxkwNPcIiZgc
M4JTbaxfs2Ecx0ounWR+FD7ARBtc2eMJJpYewR3izfYS2i4wbzLFVB0i25SvWZvIW+zVPa4WRxgD
Stgl72ZKkS+WuHuHwWzob2+vOBe99RIWlUJbE+Ykurmej8M3k7ME4j4UlC8FBWvNIu2DGr73I7fN
4F7cHeHlRMc+H4596cdJMjAEQla95xpFFTbjxtjrnHA35IQmv6WMb7QkPv8S13FWWWSpQylRmUbe
syniv4HJUxsOlw8xUeKkCEPDZ1xd20oQXINWix8FR9c9YHOZr4Y4B6+32NQApEGmmq2qGqfNvR1S
rl+vXTTVinFAHl0oP3BSv3pSnX8mbAerUN32nz4t/S6KCD4GX5x3ChongngNR1+wiRpLIVWmF3uv
X5t84v/b1x5fX3vsYGAf9OyxcSTbXVTHzI5tLuJ/EVe4kODeiRU5gxkN9KdNUcv8MHlcHBcjpGZb
G4G0tdd5Gp4FayH4frKiFfhJtumwsVoavvUstwx2Mca+POPJggcQhrjkNKe33GUY//jFwk71v/v6
FcEA48gJIhSDnbDVhv+PuH4dNcZ81P2njv7iREnH7U2VkCszcc0RpXa1q7Va+kjvn4KWsmMMoxBL
s/wFPndCiOg48JuODqCqf+2o4NyTeAkqdoSWjpZn0fVRssxGetrLxh9JJG/l9Z9bfACYyI62FwBu
CVZZPij0bllCI+Sej/XBYf2IoAbqkyMmTI/bSmuopBDnmKPR86ZN0ldQ9SG0WQzSismEBeVg2nKd
A+YcLyoFIuTzzIv8AoyuaNNPiDP7y12V80t4n3cZslbphPi/3j6RRUtP3xlEQvObS/ZkxDIb3/e4
och+ogQYTY/4A3LGHjcilV0siLQs1J017lDAt0RXtDotS+c3Ci445hHXZSPNGYkTKfptJQFKvaq/
xNKzGYLXS9YSgNerGfxELA3r1xbDqOFt9BmHTvrsIrG3dGEQ80RPhDphmWdsy1dkTFoznYxzFh5K
bIknU/Lk/9Bcco0kWl5aACqye1+nwXzPgXze0hG8nUniT5uTFY8RcwYAV99ZDvzQXTOtIkb29iDc
H0SoencIYgcoyLsy0eih0hVT7nkGNAeXHpNqGTZClta/3zM8rBBenY0BnlDokl1rVUBbSTgznK2G
WYpuFsKq/enezMkENkr+8qaejCV8hJuJnM03wJ4XHj9mzS24XkrB5IgWf2enXRqEDrSMqueMXnuF
yQnFj/eRjI69zb8I+bGNzGEvS/xm6bOGjpgFmNdBRtRHGQanURPpw7UoRpZDBq80hAbEzfVx6t1q
fc1QuxeIBQx99DoDzMcpKALYcHn/LdeinowSslz9Rvrnag4ODocdsnFj2vCu77Utchx4QbgeE/wr
jBNgKd4Pm7Ih5z1Pqr1n//Y03dne627BOT6eUtcgC464xerBmPEZewqNhPQAQ2NXpBo23cS/sHQW
/ouDzrv8ti1krQtC7tbuTQcTIfndrpIdM5a5Jt7KHbrpGG3XCKWtCHC/A66BATuLiYOU1y11Yomo
i1+mWTElXjrVVXtxpH25rcB8u+GL7mkbdj3w8uG7l3jIIeIsL9kL8ETx1GaDAdZLRaMC6Z8FeL7A
bbOLIKp8jYxFKp5Y/1hvWa+2nxB+jxKDohlW5szaLNtxK+aCXRg2Wn27eq5Quc3wmv5cc7GWWqC7
7+xTd5Le9gq+QHThgvMgEGfbK/Pe86sXE7+xS7J15oAxgNLgtI/y3t420Bbw4TNTuScGfUYHCZLq
4Bke1eJtsrGbpa23xOzKDSSj+WqI3+se6J7x7yhU8Gco+yNQ4ftFOtdwjAMkDvVnG1pLqrq24NVM
euhBxf0dwmoo0OPSlvnLOz9KT5bAv+/lW3LnF8SjXLOvcA8ljEnpAnAu4mcaC2A+1haHNN3I5Hbs
xIcjEB5cEv9oRe06tMYRchvDmr3k1GmhJPL6/x6M1FNZoa3DWCgDqwJCqSzUe4hHSeJa5yPjbr4p
4IG3FuFkBrhcKJqrXG7Ajm1Nvo/lsEdm7Sd9LbRJkcztk3pS18LkVRhJY/Pbj+u6jA0S4EGA9SQP
KOulOemoH8Cb2eugR/tP+FSYBRBJuWYyNTo0vUifzN7KP6M4v4A3ui/CPewbKCZjk9q+YvaBP3ay
ICtneY6xln4JOdX/ejWsALBezSXvs89AuUdqGhrU3wn1jLk7lzDQMmAfKnYv1ta3Z+f4O8oxSkJT
hmoM/dLt5LiTt7Zr61LCBIDmcm8GQgjQLXG3f7M6jjnfdIoVku2KgsqnfuIqkUIYRa11+0FqPsQY
C0M44uZlU3f48WAyN6XCiMLc9CCw/USrKZ1GUJlVl4Zsnmk/XUzNGsy4TYvClKCbmy0Mz6Tqrh7x
7uZSvUfoq0sSQbZtWT1YNLWZnstFCICpKM0fQvtp8xwqjb2YDzgmeF6x4pJpXtNixf0YuE96Jofq
lo4wf0b/MmKaJEHikvQHPrIIOX0Sf+BySTgnyA7UNpQ0GSRnFt0h36XwuKrwAPXwPg19fYOEqr8i
+dobmjMYg+fA+u/ZD9s8LqWRhdm51+GbL/HWLZ04ehYEhxKgflKoN2n4M/h4vKd5gXkiqc5s+T/F
lerMjPGxZIkttrND4iMrIdHc8TybuR7q5hmKRm4hWMhCaLrYNDoGAL00ClUJFeTV1NsuRS51HyoU
z53oTzTyPNb5+ONv5qunehe7dauZpqBbwO2+F2uCGxQtzdRqL7GxmVcxrvAlGIhPgIhsrrd9hmAR
Q1zxn2zPa15oNjEdr9z0R1CgPOSBynVnGyXZjM7G0wHg9UgNJIy1MX9CTVxdEPKaogVHHnms3tLa
tOQC4gFWuIl4f4JzUmUrdU5VDCfQtI3iju8qMIs+la8dvOjEYzPQWNM6r+QqjGSw1ZD8Xgycn2g0
b94mYXt0nzTyrXI87TXYXxbgH0q5vfJkA22wTrkvP88zrpUqhkbWTu4lrv1rYOK5IR2pn3N0PY1c
npxS9CkMJxpzxq6z2tYq7xZu2Jmo3kz52Z4m2RKr8veERF5/cjLRfTjqZKAsZdzC5A15JDWjrOU/
WdBp/juVrOuXBA5UB4ttubfEO1jEZm4hrMSGw2FORYrNkCRWy87VDRxCaCbhcIzs86KK4y0Hi1q1
zCz3hKzHC/cDkTPoLsAJu0cs4mkhL/yh3dqNtkxeL902Frga+fjPla1vkMGX9ojln/LOXQaDwXaq
VrJfrRlWp8bfGn4OdytOOVz9AeOC/30pK2YVOQUhuQs6A982/HPwBP+Va12oGrIkDEm77ZPIJR1T
OcuyervHMyhIMxksrA+FMTuhlWIWGCFTnKIgmFKyc6xGOvxqfxirTLfleVCUhX7k0WIt557FwAC1
atv/lfT1sOANdLdcNs2aG5VzSZjZ/j2fEVDD4AULJ7SB+kkf0oZn6SHNFmtz60OmjLDC5MrrhFgB
/2NBUVm6R82Xc4m/kUssuv2VTz8okqCVRZaA+SMsOaAgakEKYJlnit9etAl1atYtrjx/UEU38Ztu
ZCb9fpNUcuMgzLJN+TkW7haiqOpHh+wXw2SYaAJTF3SsNVi01Od76YucierhCbUf4MhWx84lNmZs
g2nLIt/xlXzCCBjadWbw4SQaSbe1Vvz8CdLLjoIGDhzz3YF47+sT1RuNI0QKuFeZHawEYoCFqCoR
mme/DkLSRrrxMKPvVK7LV+vyqUZG5nzx9stv7y/2J57r56/WcVN1mDf5uFkwPq5O8N6MsMDDqePI
ummogppDoY7QrcDohpIfVnCK3tMLFlL/+sNr5fpekGt2MP4u/ot/oWNGEikN0diWUK60cFDgJ44i
P3hXDug4DGczyGRtSjVK4boAW9Y3/7BMV5f6jRu/1btLSefH+oo+qBO4hDSrZ6vtfhpkCrSIPxEU
QkRYjVNOKbtuHZLjPjAv5XcY0juPRDs+Lcwgn7SxpAFSRMepvXx9ewPDOoWkOgNMnbBrThLpxDgA
LUXSQhvLAS3KxqcNinvqzc2gE1G/IyvhsEcY3RfWKc/xDjabkd6w4eNF0K3dRecNaHPGpTqkHQ3x
RqDQFpWe+5mYKQWot/yLp6Eb+9LRiNG8iwV8bPXiw6m94wBhScPfjf6pXYR6jrh32qDlMW8dn5R5
1cl4CyHWMGCWJ9Gmt7Wue7WZ8Tt42lBgz47sWDHVfvwj6miCmjR0LWFVubS/ulnC+ei4nc86R7PT
8AP4f/ExeWR2Jkkk6Wx3nQ+osWaHNtqb3BVufeNIgtKbh30+p8CENCzQBKdDWUsPsljmdFrhx9C0
ong++1ASBUlyC8HPsBiA9S02O/ypRMfYCyHDPqjwtgeVSQ2t8H6hNTeM0tr5K8reYUqVjnKz+Moq
vms30wbHrMaQVQq08ly+9XLOLHIQ2MUw4N7wp9t5voWFMjuAmj3/XLBVJUX5+weG2GfBS9qbTRFZ
846whCaglMkeNRo1DQ0cxC9Kxwy4Vid8XOq0PSK6n20vHQdQxoBttikcqLi40S1y9bCKPfl4okrm
+ewrEZwsG7XskEXbt6OtrSPXkHY7ZaJTdfLVt9JnusZxPQJ3cILOCBe45WILcSqH1jdeBMD5kd0B
dhByXdGzbiMrT65HKmRJLYhdGBy4T+0Hy2sbuKo7zD3Q9bBn3GfOF7FKLuASgN7zl/8PGwXBQN/6
yLSqCKx115KYnnilREhYgRIQEQHTsgYvng8f67V+6CPYxBLEZJx54a+r2YKUT4O3gnwFJgBRHtr8
5oBPBuk4MuYhmt3qTaP+bwVMjq2/8YdXsd8GNADbZJJeE9DBYpiPN4Fl2E+KcENLyYpl8R/sT9t/
YW2aML3EXv4/hQ7PrX02VtiAXsi8IPiStLtJDdu352smM9w7qyMXflA2qEn0ua4SejKbz0KdNkdg
zFAt0hSCnrJ2nK6HgqhdDtOf2dz+kAoV+yrq+gf0KbjjMJ7Hq3GuD1deXTvZLiZLSJBuS8b+1FHP
eWEnK6aMOMfYHIZoPkIREcRwjKK5z80J8IaVnQINu+eUFgySv2UPZA79NXaMNSwiTyQA5ZuuVwjs
oti2FfGBde9FWq3y2BEDSQrlqkRgMJko5SI9NwH97IdHnPmDYTFYCdS3Kvjr/KfRYW3aQJdR39xQ
1vX5ZvwQ1vbdn7nImmKLDjA+h28o7eukTJJWnxnvTeQDzepEYfTPTevLARU6//FDx1m2OktZUgt6
9RX7r6G5DRyngUA/igQTafyLF259DwjxsjABpd26PfNJ76NL0w2kU6jw+LMk3IHtmUaHuPIngSHk
dDNZG8eFeAn9/znmb5HigfE1jXjRX8E2AY7Ekvpx6J2sTwlFEAW6rmpc9WXRkapWhhzf7XscscD2
fJOKnXcw7go7lCkUieDWEjVCeObVeTdS5rHXD3YH3mcs/6oYRTu/gpOkec8iryHIiU/ZFO5qHh1/
IbPm65cCMrs5Ga3votW0YqV6DTpJbh8iUzeGa16xFWVv5Rlv5PsFeWsP89xmrDROAyHViST9n7kf
lA14NBclGa5fCtJVU20rKYfAVuQOJ+pyJXjiYBjbdnHgskncby9K5PbQdzuH0ADVxl4dmABmSxRg
TyAFAG+94s9PaYqHU24sHGq34f7IPLmYfCatznxRVeeC6ho0JAF+iLss9ZFVErDQW+UCYp6spVk2
Xd8uBrJ35WYSl0Fp5Z34yZ8TsGLPaxoX+BIpne28i9gkwG6bS3tPmUj5kd0YcvoBflTdkASdp7gl
hnPnZarx2c2Mj+W5QDV05GAIGuCTplnrWepoSB8AQncaAwF1c2hB+zY80FboQgEPuGv/ZbmCka4C
LTHgD5vyU5kdqiOyrHus4ttZuCIfsLgsZV+6wh2TJUgV794gA5tPS5Mv1ZJfcZ7iT/wH4z/y3yUj
92XoGB4tPUZLviJqHIgORi0YJQR6Ao4oc0YPc3Xh15FkTXJnK2RXGMnuUhVzPZ3hhyoflldDs9G9
t/1Me9IGjkPrzIs+u2OmO7W4PACwPsB2UbTO6HCalL6JqyR9wPjZXtxSooGf5IEuZmDyldEeFRsI
6Ec1Z3OsAP6AXouvsLPM0mHdDaTTM7r7n34NqRkYbIWhp7trEhCkzaXOikhdYYbxNilFmMmssNoH
OiYzVhXrKmSHR5MW52fagd1/eHHcBuH93miHp+b6BRz+EjXKhx9SI52nrm3u9oD/FjTXfv9u1ofP
iLoU3mrVdhbYGpy7MDq47+9mi0vzlPF8hBmlj6RLGksLXhK2PFdl+fUxOSdCWqPBNilIkxhfh51r
w5Y7nxFjlRvTR1vfXaN/91+L6uOySdmmBTpqONEJta2ic7/QbZJOYlEUplzp6P/Lq1pL1ZwQevCD
uJH00HxYgk/54i7QB0WwtFpSShapyBMFB9UAsIB3dXgN2GgM8PZl5RcqOGYHI7YxVgX+UwBqTida
qUVh1vDDLR4ax1u8Dcx3H1ZqBq1Bse0R0Zps/2+I+T8nz36Zku+uhLmFDM7MfTlMs30vINiRZfnU
eO5aFb/Jc2MZINlI/pUuuh1hJD2zOLULEZXIsqPKVDBo3VSbhyC4Vrq2sKNer34i0vAR4cPloAtX
V++Ckm0BSaHtGf+v8y+DzMlY1vYqMsNUIyd3o2LGABUocN2+OJOANuUMcV0b5wy9ymEk3fYjquQU
jlnHlRTx/UGjCUchZjByEFDq4ix+7YzoM0yalyZ/hq/UmdHe1ZzS2gxjdYdqsuVMbKZ/9U/K9J/+
3DNAS+/ObX1VFS1EckQI8J9V8fCij7sEI9H/hH7nRYnVaNUMBdADX2ISBdZ7+oMkO98eBDEXm1/n
fRZd4TYnZOCuUeDehZQKuJ1nGzNIbGpFgwyo83Q9WvME3Xmg3sLUftTwtCkF77VB+YFJOOv+Q770
PCnmaahn0KEjLa4pyXp4RimEAt5AQmrXuxbZuc8q2Wb+29c7vgzlVFbnFtZMzNdgIMhBBwMQseFY
x+t0gMQgvp2zQwTnCWaUeH6M37fmpu4TjrWa8R/XTU4qWcJ++zBfYkSZPREH9GuneAaFLZuYJxuZ
W2h3EKSZl0dYAkV7OMbLLAprRt7inWs/Tcv8cspTk2RrXmQ79KoSTN1Sw9rWUdEJxJvwMiFtwIho
5u9PI2DMMYhT4GHIjgoGS9UtHkc5r7GB5GSaEtbASS6irU23DZUt/YRtRdOrOIXwraPHwjPcVIWM
hYxGuJSWPq1bDpeIDI5yaj2Vs39oVGWQrF0wY5QpaPNgld3uIlzYJn0WtAhhzOmFUPXzOcjZagZo
aCzVYvvX++rPXcZJmskVP0GzibGKSCvzSIy3HhV/9g5600pglNvO6tXQ3zNWlwkW98cvhcNj305O
wd7XW8Eh7cUAStTpaFdOXtLuK47R1qEvWxwrqKSR1RKjaLz2JaTuqX+ojooDLB6vu6Uinuo++j8m
NcLxUlKMYeLZpxbKpa4bpkbUoyUdcG4Nw/sPjzVRX2BG4jRSGoA6MonGHCgeOOX/jxrTQVoUiwA5
tH55DCpOy+z4AZmw/4IspAthXtP3y5DbIzH587PBZlp/mblktiIWhcTnyJeDLu6tZp/KWYhe9Yxh
48EqE2TPNBHmaEW9kFKh6CecNyvbslHnG7qDQErwgSMMgzCv2/w5WhWDiKHiwXQiWAu+PEfBHjZZ
/Z5j0QoiHw+1xW4W2XsGB+ccW034EihiI39FvRnmogbQmge5tiDWIgaEOya879nYiBOYN5UYur0y
U9fc1dUosAWmT3umwaqyxHtVYfPrND66Wb3yaauTJs65u7rdSsFGTp0FRqtzaM5ZPcANAUWzfHLH
vIQtOsyAFmPvRgWweaR7wbVpNK11lZdIxXKoXby6uakVaN5sX5zXsg5kCvnZefTA+rnBSWq6ZYyG
2wBSpR/eIcJxGIUmd1Ma5cRRgFT6knYmbO93l/GShUjE9H2PAXtGQyl5cYmQ7khDXJK4oJlPs1h+
HFxiO0jjI1MeqBlaB644iEBs4x8zmES1+zJ5qNA5upSk5G+k5rcy0+Vm6+o1yXV3C2P1geooJ0qG
8aaUZPPX+/cfBh7XSNqe2mApUkihv80NkPPjkja1i94OA4ACmkLq4Gl5Miml5TyC2XXysxevpT39
iMirYX5KRrqvuuDxZmBdmyQ3GFZLNtAt/TLGmJrhTi/yi2C5NZ0fugxtK0wb0EHZwMVnBdg1AvWI
uydv801Z2iSY6ot6F7+QEZfZwt7J6nc2MyiURbY1G8TA/UXfEQ6+KXcm9tBypid7ftJAfhG8x1C1
/XdXKy1IDZEgN2CEGoi0jYNw3lYRV3+So73pQygcKMddDSgBiWuiKvYXcBdHK45agz0rMuT9akcu
PYn4cEjviD7vvp8Hbx3Si5+7eTckTEAsieHpVB5eFpLYJIllqIbn0mguYPUWqLOZG8LdvYySp3H6
RUMJMa3b3sQPVdnkNA7BlYkV4eU64ive3JTMFq7evTRwj4ikWyh7qKlNbCRrYjek/WieVTM22wjW
9qEyNfkOfPglD99s0UdOuorfIK0wlNwJlqEBf7SH19IIfalM700UUBZH7nyPXXIyZcaDt54KWHLf
PW/+Pogj64ikGxmAEN9Ej4ANXcNZxQLn4A4IgWW+rQuKOmzBWR0IefKYgmcFsNVaPyBVXpMSdZ7Y
SIS/xbmiB4p2IbU7nzC+BvyCMMG68qG50IgiXK/tjDIHqe7MKsh671L6x+vtB+oRzUA07PpxYLIK
NcqmAogePt+5XBcWDP2ZPN86moUG5psXhadA3WyWUx8TXdB2if1xbGjFQPtp9/I3WewaHZsObUHC
3rF192Cq5funZ3xDyAVizrkmwgwqwvH4QYohdmCGZN1X3b4H66Wi6CwI/QZgiKb+0heZZbkJmCDC
SHO7sxlJRcE7zKtx6keCte390mLwS381XzZ4/w4JppQImx26Fie/EEzpDvne/zRVqmqn+za5VSOA
z13MtWcxokkv0guc1+dqgDFS9EOVPjSqhSjEHH4rreZAH6s2Ao8EqGeXAbjf+oAvYXhqhutuSiTj
pyWK+FRsRE6YxaqEj6XdmHO28rh1J1W03khkkFNeBOdhNXtYj8gmrGI8URtVZX3Hjv7VlRXvKfOB
56CRd0jOkZCErbgF0Tm0C5XaFBeLoq7Cw+ihV5mfRAsGsbg96wt8OLBF+W5MeNpp2s/RTj3Jt01h
T5vfqwhp9Ka5EUTs/D9mpoKvxEe6WKa5YgpPl5qN6pZ5M2tcJTXrHVTgAV+A9C0z0j0LuDT4DUbF
W8ZnwuPxUR+DNeQmUrNdisiFlX2KuX+/YF4rIWrGaEk34vbHP7drpP73JKqG9n38rZaKjOgfzi+G
vOpj3pDoD75GUO7ZnRWrwuBMzopNS58WewDtZekvZjaP+2YfXZy2L++J1nQfpLjMS/7790yjJC0o
MGOtYxg1G4e7cYtAZfZhR2EOP5yzTzOPVpdNSOESqiSNX/IOktvmMk2h35T8vgOtWlhYYRDOZci6
mSKcdZTurZ1DTf+2ZOS5UnUn5fRZ9vrbdeRv9Yls4EycPUuT5L1bIXQP+MnvtxT3ucALzme0dOZT
kBrGmmdnNFd1DC0K9kE4BWR+XlU63asTxwCgDjn9ZtQvQ7rMk3Zj5Vfr1DoXv4Ylj05+f4hNxee5
5NQyDhSwHgtlDv0Kd6e7ojp1X8vouhph4yyJDc/BTtNig1q0iCaYOi9q7OWN56rYvi9PPbcLhGjs
wvSVe0ZZ6BfS8jEUMnRa5Upj92jOSJ5PHXp5acNT2H0vXlyQhPkghdwEoPNDWsyDsqgbXv/EorRZ
qiQCyODu1bdCogLsVFCTdyiQsJ+fRPIzi0mEdQl23aEVRyRinZv1Mu8aOvWDee8P37rqXb3D6nE6
abvBjLCfwzav1GqW2yiRFbR4D+10gc1CDISjHWuJgP14MbWQC8T2yMoVCUf1S2PL4Dx3Sytebd/I
vx6jifQwRA5+gAZJNTqjAhyZhePF0tfrrV0JJCSWDE3JD0kqgF/PdOLp7XGTDI0mgzqzX6LjH13K
QS9qZyoA9c8S8nATJMltVQ2cSP8/0Kl//eB4YkSXFhfph73yFtckAuVB1D5hfqSc8GoT77Dr7k8l
G/LJupBbZ2oIy2TVUbMR/1pYb8RTevxXI2nxoz8E/ahK518AnHaukJaAoxs1KAxsWWU4upwrlAVs
v9SviM0wp5OxTXfZoNJelME2w7kf8HhY0uCCppHN5mw0Z95dWkuhXOUAdaueba3LyguwNCS9W2Af
E44pj17ihJm6+WKcTLtaG8bhjCUaAywjCjdgovx60FwdOkdOBu4BihozzUHjSfC5/grNuFjLV07E
waXd5TwBrnnDLuMUKNPTmr3SJkgVIeobjIn7I58e7PssS0T5bShkr0KJUENbsBeSWX71sw2Xnqif
wqwemkbvE7TJ7e/NNe7Gw1LvD9LsXE3Y/4WLML5O5ngAUqOMPX+FLI+RHqU7SsvMLGd3ehsv4pS3
ESxyh8Y/bBGce8PJ39UPVLOFOS6EF8IXgeKZTTmOWa1aft05UmpO7j0fYsTqIhW2K+W0Rbyb6ptd
iijp6LZd/OzhRzLbppwiSt4XCqJIfNRERtEAlLFEtGsYWMt1yn7lvCnezGfpZbunCCH8ea1D3myI
WzLf7tU8ywagkmOMzy7Wds5jssqJr+6nDL0zO3ZYH29lt+JpaXZVqo6lseTc4MgerBTIWbcj/7rP
GKsMqE3uuv2Gz9tbrsJyqAlbWZ9lXXmhoUb5J6E/XoxiqnmtZ0nRLgVLVt9v0FR5zDn4S2yPVeoA
ylFGZWNboDeV33S/xMg/2q8sIHYUOt+S73bYTougO2lsQo5pdIEuEIQODiX86B0ELuz6FAdlwsxM
ZxzQp2WQgkjUBuLgKuXfzSCBjZdY6yZfFrHFmY3LJYjSKcW7TcjjzrgBX7iERUKunohhSrLmvIDj
X3lH+Wj4Tw0V/en6tUBcczYJUp43ATfmnW/aXaRxadYrK3uruEr/RPkamwTEEM38yQcUmSNHiX7G
o7/or/9JM/QNZLv+oXpkxq2ZkDu+xzDzjPrc9OThbKKjKpdW3gPezbgNl6F4drBizzDk2SNWD+iE
VXNK2WJ+2On+xHxlo5F1M2Ly4/ZrqrzeZeJCI/m1PkDA6geqq0aj8oqF7rDlpkrOvr/jnUkCB8bx
e0RhpAKcbLPhKE+tAwItfzxnpK5+TknX7iq9TI9rjYBH8NAmlHIwJvf44RpEAf2V4DFaX3V9dPRg
fI1LpJJqiEREjOb9y50Bewer+5Mg5CMjiUz7DLW5p48Io6RpAun6QW4bJFQ0NETlbEdJPNlCiCIM
N1UhOOpuKQFELyoEVIobKeCrXZB0bNN4/t1d7p1y726MbhbKIL/bQAEZ+cMOYmaaut57Ksui+Rxj
17y+QsZQBBAbmgZvnhjy1NTP1rDVg/sa0DCBH7k=
`protect end_protected
