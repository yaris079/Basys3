`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
oT0z31FkRWBnvw8tQSYlPgvwMzQiXtg0HPkxPs89zOg60hrmX6daaxUTvDubfRdFMPUqxiU7VqWR
fOz2cmTQkg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jO03cSr1nREj7MKe1Ki2/yRdN7u4X5FG+MPaJkHEV/JaCCTTqU1ZxA6HpCI88nbM/S7h+SvJsbPh
IZEe4btSQGTH3MXDqfZAVoRuHikRAjhkufFdgp/Gdz1aauMyqTCNqs70lZsHNNNzkZv4GAicyYyo
An3E4KIkdfoCOXp8tFM=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VOEAUxGbB7UoRGVW3zm/mvfW3nULx1THQ+tBcTOEXjMTJz9IZZgoTGRVhd2dUAFVqbP4Hog9wJNE
ta1m4ZH4pFiIHZPdq1H5spGbPHoHisJpraJqBd7BRAUX8Go2UO+N7r50QsjWYT2JE42jHVESAJtZ
FCEM3EwuNchYSHTmtET0Yzsjsx/7COJUxijQS5BpWPZa8eNTJere5eRcUjOG9l1QmTO8cxA1Xb91
kfwlYXNNwaWvkDHDvHXSyv8yLV9k4SBkail8Op0Of29Eg4nCQHqCyEze0BzeWXkEokRTkINMWk1k
YHEPYBJLTiKnnR/JasPyCoCG053+UdiyZCBlGw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2hbt7aoPR4vBV7PsDyE4OLrVCmNJjL1FbxJe1CtQLmuOPole3nCCRnhyi0Jb5/RpeSjuIygaAGSa
P4PhHEChrH7ajnB0Ze2+ZEj8NMWF4CjC8slEWzgX6W4Ri8wZf9EBOnc91ikQSHlMcEqdCjFtx//c
MtikM8/x+SmxgmlfR38=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YL+q66BrJK8tI6jHDJmd03rIvs1CGNbQanhCYkSOcGqshSvW85aueeQjVzM2/ggcphtntpyhxnHx
CedWePZjAChxTbzmMFX6w53W7MydDNFpcUa22zqw43PPQ5PqzlD3v/JH/EA3GWR3cqjIPhXcwLP/
ZEVWI6VhMeRzuMgQcz0jEvP11xCf4ILtPJmRCoT5qEpdOdtSUlOSLr8cOC0UTjmQrZEipTtwx7jU
IAEo4N3hLOmezvoUEAObWBgAPzDIF5lD4QJHljFNDlkQ42mSaZzh+eDaCp9dCG0QO4hIIKcu93s9
aFwCzR5z/iLiFJqEN/OTaeCv5UeXPQMZeMJ+0g==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9104)
`protect data_block
hK5VRKSatmua+so0S2nAZtk8FkcD8jzRoq4+2XPCWChnXsVOxYXFJAZdcqYhLmHj/mNRzXu0lGzd
i8gLg7o3t8dsoUNQGGkJDW6pkEJLBkjxtvQrLpsqIP/nAHrt7u8VSLzkV3WsaPiZDZm7OK4HUHzU
FI245PqXluRHruEDpvy9H2947gvAxgnVpoTz605ERcf13jUMUS1VGFhn5OSXoc87TshTgDhk+hw7
bmWMEe3nPRuzhv+DmgTyvF30ijCbJG/WbseZyUfNdGqVI+XJZaFZ5z+bVGhqD6jraE2soGXKKT3L
7g9BhKUE+Y8VZpw7Pr4mF/ILxiYUw6Ton52RXcmuyE5vBhSq/rfOwa/jnZC2ZGv2cPKRuVHd/GGD
FetM9u5HS1jbFhzhMn619e9zUpBk4iy52a/JIjdstbznYd6/63mqRzpb2XZJ5ZMmM0a0C0Wo4TYe
9hLmfchQePtCMubS4DjoOHoV5oqH15RhcxnrPw9QiVMGwSzFrNRLc9vQJSa5+18MkClNeOmX7B5H
BcAhs7wzKyd/O/nY97P8rOdSoYUiAbsEtrzsM0TmTOezBcA5dnqAUoo0b6M8RhikQ+Q7rkmUCEQD
hxANS3vT05A3wFriWlqBfoVPaZ73ELPcfo2mUVz7wMk7BjJ3D8tY0h5rOy3PamoHofEh77o7DxO8
sWk08J8F9YCf2buvIQfzvZRWGUhjTn21v6JWgwvaLuMYI7F/MrA3bz+uF5aCdAvSOuAKZzfr43+E
n7IErIXKVFZToAa92Cmcrhbgb4sIqYPJ7nOBI73ky2cJN42CEacG2Z/a8HZoS6w1ueF7wGANLYmq
dzR1X2wrXjhJCkBNTAeDYCJY339XKnIJNifDFTprNS3jgfG7m/ileOEl92Wmei1j1mqmcc26pqR2
/G/uwq8VB9iKN5ncWvn5gEkgMElawToS8uCctDczQFhBlSZSr5mGMawho079tBHy/kf0Bi6B+j7K
NkO6kjKXQAcMDtpoGdDy06/cDYArMzHNVbyotATfsgMKk/VorNOPsURVadIydv19hmsjVfZaxtox
sVktqtuVkmgewBqYFmq0ZsGi/NmRhZ7Al3m/t3JLxbqa1HT3ytTi1DAW95gogbMXqMuYgeHSBWFc
nnNX5hJuAI/NP+pJ07LrGrK/D6bg4KOO9qp8kWyK3CotaihpphLcjns0LdPW7VjlyiAHqtoUZXo7
BEeHpGZhtphjeRw5bsbyafePBAxaXLujdunJrI7oTRPnSNfNy6JSZTomzuDeUbwwe7m9oMKunEoy
6ifOgyI8JOvcB38X4hgKpUQlXG7wNjJaQnVBEs3tfg57pof/iqfBXpkXeZxlLe89nOihJ+Qj8O+B
0wivw+4w2ipdHarTUVHP8IJ3L0RQpGugXXIH3CitSxqwfe1ULM1cXTfbcu1qIk6HT03YHWGbYs3x
PLjHlhU//QSm0qP8KPoZdzI8+tX8ugHMlNkCVqb0nfGCep8VuYQiHF2HNS/LAy6qeFNdHIZ47Zn6
zREhA4XpZKYYkKtcE4yv47G3XU3SFkymynI68sOCHuD4LXkN9p0nKBXNf+CZohgMvZ6AMfmclB0+
GWJi34dawJtZ79MItF7Dhe53bW6+a9HzVY2az/tWBnXnidNv+uNgCmhG4t6ruzVXfsXRoy5/HMKD
dXwOwraNRQED+MT+/x8TueAzr6IE5OLl0GkBGWWyCBA/Q03Rl7AClHilrcwsgJf1GcIWDPC/fCmh
9dssiVWHZ0NVPtZHsPsS/TH/2DkmJN2MTstgDx+UnjtBJ8tmyvULEr8p8JlIAOcPdM6KyzDKl6O1
0CXoOHpkWy4cvb4pux+AweFJakxtX0s/lVVZKkdxZQ6009BeHEUcjK7dki/EN4otqDaahCDXGZTA
zpFcywK7Ncmrw67ku+6sygGCT6j7F3tNjMntdH7GAXjPA3NsT/pnzKhjoHc9W5GCxFReV3fs3sro
AbGAfF3NbtxNkkrmrKWEjKwCmFzZblRBkBrjmiqwe5joWtAkoBnwAFLqspO7/Z3wPz8Ujwnb48Wq
f4qVNMvvqzc+JQwgkoWIsmPTvyyZXDUXFJc2Dqg6GPGoTAUFFx87WKlZZL+irmTbWnmq/t+k3YOm
lSq5OKG3cwIckBYXBinWO78Y/ZyaTG1mSzZqk2zRy0zmfPo7rXkCvzzZHopMJKOmvfz9sE8bibsi
4p393kw7LA45EQ4AWgpR6wv4eYKSUrEPD2k+EWecDB7UC9U6vxfQBsBKZX2q/5EUZCVYfftjDEZB
dx+15kmiJdplwP6fzqbVvkqS4juAmqUHcu5LeWOVNDQh4bNskf2IFuq41qxdSyC+q7u40BGsqP1o
dRDUak26boHozIdJZvH2sgxa2DJkrt1QEhMrZoMzx4IXkSqnqzPwVSxZF4MZ285Usi14Z65POUbK
sUL2PE5kugkJ38KksdtlMvjWjdDXYzHg4RsX5mBnirHo8H831em1AgRd+W+gDeF3Y6HdfNd8pbWz
mZRYfKA+slouByatQmykWb1kU6wxL7waMoUEhTHjfW3BvsHvZCe1p1htsz+gmSfDvo0oUQEmqFS4
Gcq0AnU+6YV5ZmPbmuJxSz4TQlPbi92YxGc/O3PYVAXvhaCQf6jDwJIxIjeMqSkG99aN83xKAz85
ZRNvufI+svAxBlVrDPMbAWTSdlb+91PJmZxRLSa53rnO3QoUf9mshEkppfCGl8mYUhX1YHHauHO6
d5BNxp1BnkXnp3zYakGXiwVR7TNRh0HeC0aC4mbZXSBr+YuwP5lgJ3woNLR/XJhVMuGqp0BVVA1r
jIcIxBjXCkKpEgZ4AZReMxsY6mITSSVSYtaXCdiLIsyNyCWa3WAkUr94RApyg2XDKWFBd5hhTYQn
NiAFCDZAjoFSPBTzPpnzuOaPWKwFZOFmRX9ZV0uxkqrh6t21o02Mgdv4EEBCTXKY2SlIGwy4f9RV
920bcPQCVe9dYRGysZMY9pdDoRozA4RseydcU1dEhTlckWe06a42/dhm0ggrI7F9A+zaSC9tGcqJ
KQ3GNnNUGF+r2bgBWTSkp9KYWz9ziSYQd3SqG+KHjizBE8w4sdyxcMFOL5T7Qi3G9WnL/riKBrW4
2IuQSrkIE9XUjlq87OksLivgCQ6Om/VzJWROfiTF571d96SGXsScGgP519dkWmCdC7oImjmx6KFD
PKG9DyU7N3BN+7CzKqIykKJ4huK1Fvu+Rm0gALfERYIVoJ0jqYogEoMqvjWWyF14CAUrbzFJ6AG0
Vd1+rGbJGPU5v+YM6vrWpp00Ws7844mlhwSNAho76gFL09J6JkZB9n8G873bU5G0p5pCWFS5FmK5
ZRFQMzY3+8ybelZ0YaZy/7YpD6U1Kff289ReCz9iG1O+niXc9p3SUWT1IX/+dBMgPYlu9gCGi9m/
aUi+Z+0KDP8qCe5Vjkt5K2R5eXu3ycIyDM4WJLu36pvqi8E51IBQCJXGgH39a+wkplm2t1lONnA9
hJLgp0dYJEQ4TRoiP4JtEfNxrL2ZPUUZ1VvOZIg7rmxMDG7qoZ3oI45ihZOQFYFblG+KIUI2Dp1B
//HdMdKY8XjZkzuJKQDgX+kkMiN3316EBGFmd8Be+Ni5IJwPwTMOKcUfHnC3Xy8RHW5nphJDZMKL
zO5akHyNn+ebVdu4JWH9510IMVjUqmEMntmqY30ueLADPR7tlfvxMv1ezGb1Ktu3OGgHy7A15B5a
5th8H/jClfjh2UZXos3wlBlCf5QZnU1tDfaBpsY6S8ULS6pJqHJzVnRoQcuo64ZZQQakrXim13Qz
GVl+zNB4eBhuEgvjYIAudb7u9TtlzCD5zmcP03bhIZxbIqUMFmHjmtmTDLKYGpzwtxVK+xVcm+a/
dXOcZ0ykbrAIsPnyZ+p8moEGn+a/Arw6CL0ddS4v1jmoiOlqMQa2w131O6zU8ar3PvAnjv/TqnB+
0x9caauCI2V39b0FXj+xM7LwK6hLv+Se3Vd+aonPHfQhCIBdhWnUDtkMDoSVBxxba+k+KSQpTXE2
LPdzZqHMzwI+VnInlJGzRfHY+Uqrqk47kSEQcpJpmTz1WUP4eEVhohMOmvHT7/Q662juBY871FRC
YhiKe1x3qSgezlNk5CobYX9QA7BP3tSSq/DJyg1gA1tSaVtAmPpTAwmGus+JZsmCS8Bc/4ydCBL/
8Cn2FeSfQhKb1k8bIHJWCaKlwOUOR1tauoQIiTDrrJ/7kbDdhfbm7PAnIUmmqsypdrS1hzA8UV1s
vxAeLdF2D/B8xMzj+PkNHgZnwuPSnKfgu+4VrCaS0hojMX9RBcIFIQjMkRRkiARunked40Pj3rVk
QVfRPUfZFaCjHu/LctKQgjxu5y74f1UMTZ7+W+brIAjSDl61W3HGQuvcObJpDtpN8pxlctxjw9vl
wXfJfdv+nucf6DqeealSSsEBc5YbVlajlF8LnzrBgHks0GJsH0poeoXOGfFGA27wHsovqnoR88yR
/8YfI4KBGNMxLYBNtv4oArvNus9X7H2U8kETiwqZgvhF0FZGITO6ObVnTHRLnvrsXoquwOzI3HRC
l1Yv0Le/rNJm3XX8FJ4Z0HbgEe034jorg0BQ4CZZKnFcOPmwNAJrJ19/a3lLxbEHO+0/s9cLDcCx
YyQ6cgza5PZUYABXhXPfPLR14X1Vc7s0xTbTsGaWRI7u8QAm5AJQNcl0o/FIDinivl/uC5J+CPBb
iu1hRX3+BvmbYuzxhET/d8axhSrilBpyPsfVo/5ESKHJY0B54kBFaTWG00Cq2GL0Eph1buIFb/8b
QO061IN/qAQrJn6x64wJsZWh6BkoJth+KHp1ViU4QoR/JdXnCkj2FIHOGc/TmJWTDCp36EgNr45d
L9WyM2+rO7vJBiZS94wnAcJCPhrW18YVMqCL7JQET2/Kxvs57sDX7hzEuRJW+GYPjWpPjP3qEG4K
8dar8i2377KzDOLRarlllsTUTtCM7ZcJFlv7s2KYZPk6YC2OUOXMWaFxnJa4En/oBHaNxGztJorh
X+uFO4JhM3O8w0n6bCjbK+63E6er1DDP/3VcSforFe2waZnzpcHKbhZ/Gn7T1ZC0sfGzDUdk7qNL
1Daag2x+0lWXlkJ3dA3Ev31hVpcWLPmklzPvJw3a8I0IOjoXzg7aJm0uppgi6Soq+p8N5eXfcl19
l5yV2wrf4XTPxsbPGYzgdtiU7XDaTcU4ZnIoG5qLU7otaNjXf4/Kt5B/x6w3/vDnNVhpEc2LKjnk
r4vOmwW7Hx8D+100HqACaXcla7GEA0AgV5wl2HJq+03SWRzB8D+Ht93bHTE0EI4fXmzgjlRFeFIj
6LwpMH6GBxUbWBU+rtln8TpNWviCkl/HXwqIFRbzdbxGLQAjkoCKy8q/UbQaxnfcq/w4mlDlPEmN
KiOeC04+B+crtgDMeBt8db71A6jL/iYE8ppAIiX9EyOliOJmhEkPTo9ce76T/9rB4VnlEOhUWb/P
/Su4DUAwzYTY5q97z4L3SmYlxN2RXN+0hv99fFq94XmQPuojQ1W4pNZtA0GOReE04iNSyrNetj5/
NDfeFe7qUmp1vSamKNjgM7pvdsuwiILtMxwvSYRk2TUmF9at+ijCrFYMVhhWm6fJ61qYztxNl09+
CDFhqOr3o6j/psufEss+uUmhgVKx6Z6bodGeInqw3QE8sTNZ/Yejph9NotMHxD7nBbOm+EJJ/lMv
NuR5jkdOLWrmE8Hz8UaK9hyQUY4bnIvs3OL0DL6h6BcXQjc3CsDmnMDYAsYfGvUW8NqNlPWXAfO7
Y8OujFDvklJrPShEf0gSPy2KsnyW5Iaq2HhKcGNGKwzrjAhTDt7s1ovSFnzREQLYTJbtSnsdV6D4
jTdXX/RynIzCxwtUq8wADftVKFy23EihWrPwM6vKGvNTwFvXE0wpYyRkn0SMSj43snwI67rbL7+O
6NrE+3DaOhfYWuZn9iaTy06nJk5MVyJNuKvZ8ttfJKX8CLH/Fni8HrmdVFlgSbd+Jlp9+K6uF5va
TPjhuY6WLBogYy3CD3ksgGC6WCK+Q4rDXKPDW1S4vpaR1CEV58w6l7zOwhxfKJSFbFeCr/xNnh7z
dR3fCgq1pCS5sdjZ2vGqbUoupu7UupAJRMJGY6bmO0d619vfSr12r+QAl+Lzf3b7v+0dREVLMqww
q6aOI6U8ISYfjfd8xQkAZqjF0MtSh0wLd3Cd0rjzfjJ3p/+hw+/bPyJHD3Mf1H6SVpxJdOkUt0ZS
gzKwubozeCush3Mo/P9qCpLSUEDEMj/RJxiZFQLlu/r9haU82DVCWc7RpvbBQoMH8ZsPyFrGTUZy
NkHVG2bZpJFD1A5icRxYjBtX5M4F+dxllq9W5B7BvZXNIFVQLFeTNhC6abCvvNEttERaV8cTa9kC
qtpxlbcC33/qjIbAvNHLHrq7UBT4pWfnpwomutFxYmBn83JrMu+zx9brr04IWuBJj3QeW9ZyBJvY
7REDEUXsPrs58NA94wJ+PP9T2WvTGFhcYX0SkzWkPsbvxH0nfB3llBsP08GPvI746m6z6xeU5M9S
pf2kCx3FSNb8Du8IXMIwgtEuD9Tfz+S9OnX8eLh236Kq857pbCEeaq95/+cIE7nn+kU2QIeyiDpY
3QX4gGxYzb4LdMzcLJ8kVF31PkqeoW4t6fKjdxMEMZGs78sX+ffcnw5yUkj/u46TycTQ57I4Bk3D
SurBAWi7jEjQdR9J6Tl+j0Nyri01mtCtfXNEelfGSqqr0Imj/d0rBI7hBZdwbL5EM/yVN+0m7g/A
KmjpVUZwF4+0z/huSSnw439+fdI0/RlwWLaDN/8RE086PKaHOglEy+FCNnfutfi5UpISGgFyPrsx
X4N3pU2Gx4mSZaorA/Q8WONm7FFz+oJuzCokWRnH06jffwJJUryEB/OlReDr4OTEAtQN+exlwSvC
idCGbAeyOaHro+EGS9TxSt3y/tU26TFNrqZzX8YzxFa0HMiUK5SCtprDjVkAulH+5nJBksvpN5Gn
y0un+4yexQ8Kkz7QaFPkhL57z/JQJHxmyyAH9wMWhyKa4BlvQ//BaqbIe8umTgQs5HugVvQtiOdm
yAXRHNgtEn0q0FA81oAaZCnrWoPLogJB1YNwDCHdjHCqTMvcQACrzOG6zZxQru8Wd1xftYV0EBd0
LhzAniV1cYjYtZuZBk2/LTwqWv0D4mVtMTYquSYbvjbSUuyeY25nb5jV4PXVvowsYDs31JUCAVfs
nzd19i96LxFlLdDcHkzwoMKBW/oEAEiXAhsImQOjhrXezgRtl2AHqT5RRUVHTrrfSwCWkxoYw7i8
Y14msd2VHSsi9yHfI9zC7yBcMT1mSOQgI9YB5U2pHW6Xj5RTikRf/5RWdDOKciOkB8Rskf+pQaSd
anOc+WXyh+lfWILAJimCk7NukZQMfvaKHOLMsveKKO4WV3XoA609hSMvFmPe0EaD8f9lzfwYy4uE
3gd6yeN90w392jflHAqL6xNa41kBqJmMwgo2CVHhm0P74UfDmjVdRNfNi/EcvT9xbHz77ZYcsZ04
23BkoUAMde0WnAU3H1eBhk8Pvb9BeH1uMBuHAUgGMrAvXI7euKLYWUBdR7wg9fCdIaQ/PSxNfpRZ
iH4TrcnorZGFEbTJmgYADM6D3045sBuI11RgzsUM49YIGXf15guqR9V1RLlXFuZVO4ENE28AH7N2
6NATsKxY785kX8o6W4CkDS/zzx3UQiXjrJkSQ7o7eYbIx+zT/uvr7Mo5lndFDrh313yE8l8IgPDj
KFlawvKZtRh4Z1ECzH0dVbYaj97Oivu3uQY93yM4O1csJmZFeEaZpFcczJnUAhSezV2njOQEraVJ
i8lASkxEg90KnbEhmFD0bQJOgZuRk9GCwezOOHI/th0nvlM3o0j0XeBFbGsHxfOtsoiicjmp7igf
0X5+AWWYtz/dxREh/DeshJFNSaS3iAgu+H26X9tL0mCwlI2/PCaHnb+QkYLQjMQDbHOBggaoSrAt
xiL8KDHZWwg0hgaN+mR6QUHfkgEPUhRV502cei0lDA9h/+M/KXSgLjkSM2/Qd7wRDMLbknQNHXc5
yonJN/HYAz3gqyLuteUJhNqEXXAv8YbRF7Gtlaobm39Eq5EIJdaTofOGYyzVPXsEbA1lK6L+q9bg
5IFniz1jKBU1HQ5cTQgW0hWIYAIaqoxLl7LPpYTGEz5mVFTt1bn7OB1JUVAfvow06ZJbR4uKdoQv
AfNolBLKhmlkTqrIEnwfy+7qJdOMW12RQC4+e2cHii4sgPcQ8nzwfGZq5XBHfVj9PSTbDRXekxnU
Jxwg/2V18H2rP8kraljrTB0iodveBwkBnG1crnM/8/zle91uvycessf0moHYR567kIigTEtMJnDD
A7FrEZRTgLu81Lrk8siCts7ToKKVWm/M6YZB8IrlTlyErv63Vy9+3OvGSoh4IYDe3h/OFD4L3zkf
zNj+sCd76IF+GkiaPAhWsJ5jdfBG2/JUeTPPwzb/VBpc+O8VIP/2itVFrA7TVh2DBzCm/iJHaiWa
QpSpBeyFaBsQo4gorQegPTFqGaRa2hwGF7LHg+oHNUwwf+a54xlysQMdKYQeIZ8gu8EF/aCnMfws
0m3BVq1DCvgOSv3lxf/JH/O+LefIDnMu+LQJOI4CAXWI3DEdw03pQXR9dHAS13s21CUUX5aHuvR9
vs3NPJcUSvR9pAe2MWoyrbOBgscalpNz2g83TF1C0R8UYEWiclOvqva2p/1ysmSk3Gb/pw4E6hsV
WVC8OraBWWQzm7YLrWujAVqWe5dFYakI3L6AeW+QbGi5r2KehibrYDc7kKgZEv0R3YLQYIV035kv
yXKbNDLAlaQUyz36KItwqE1zn4Id0GO6OSQc58P+eOlgUY8idiDGreg/mYuiJE+aK3K7akx1gOyU
c693xHPW2FCGmnvdhQzJtbh48mvQryFBbhXWgDB+kKdnn7nSPZKNppNzs1W+2YyaqtE/C59vaHyW
1SMBB3uhTs28d0g2HzG7x39iO0rSBRqS+RWXMwsU69m7I0munm6jwwbH00A2xKX+A+5U00c4OIzW
417+sgK7AacY8Z+TXgYylgt/0hgf2ZGE/8kf9MKZloCMfxCccFfCMcSEVX20cgL1CEJ7raoDs4WE
6SowZp0cV+72ayx+OKHJj/NMgpVKP7VB8X/V9ZRPTPDf/Gq5AY3a/p1BNLdnq74FwJsgVPFJbVRN
EZa4xFFUfkwhu/BIxLjPDnSM17lYzyZvJeBAuKoyQJc2+QBi2YV8k/L5EhK3gwqQX5F8pKlK7cfJ
hc+VXNJUHLLUFwTphFOn+Qx7O9HM7JhJz8ZhXL+r4Ei44FT9JvvYfGUuyvIOT5WamzgaBTdTE7il
InNlCQbt0sDh0DIEZFywZ8ngBKc2txMQTQfxwV1LN1JPb8lZgIR2wpLQVlqOkNo86HRkz3lBBjEC
lpReCA2vU1uXg95KF0imm1Cvib1noYsWyeW139R/AUpPsBWzq4Z/zbH2vRDCW3FGKTKo1xNLEvt0
RSiyblHoNyu+fzmFCGmvqM6GEhAH32ThsTMwMAkSVZ94eS70lePGlcr0GD+hvjVEZEUJM8jS1XXT
xdjk6pquIowWgsabrALUbvrWQ2GLpIfr2komnXxl009n6Nx+YsEIm93TCrmcnKGXIoxssttC9yYA
ssodiRnreHO0Kw3rND1FTyITEdzomU97gofh77h6DT9+zB/qH6kMGBuM7gR8vAsd5mj35nssfx4V
Kg1XrzR0g4qVOPiWnhEEKIJZAx64ockcpZTwkaHop1BYsoljexW7fMziLCNsTt6/K8JVnClQdzWu
AYBrUUZbuTNWX8fh7hLuDhTzFM+JufANoXFoMxwAQmBLo9vcT7p4kix6Gyhi/xYk7xdvYIzc1tL4
qLmTxC/KWjM8jyWTq/ZaH4YD8pTR5jep7Nokro1bHbkX+giEPDg6QMBzvgO98zQKhtjyjjX0XCS+
wRrga2ytuTFKqQg09pOg75KIIboUYV6NziDgqak3Sz0M4C3fbjLRIu1vrB8ma1acWKsLFhsEdSck
JlNXR+9E/GnkEglkqTt09a0owGDnI5jHm0OiruRGx+E7+GJKiBhhCGQnMtS+CiIje5sLVmPPLwEv
6I+sUkvMt4nT6SAxRBLP5JSrv2tdM9DVf4Oi2WDBkcJwijsKt7pijVnOi3z2W7nb9q9th+j3h8VB
QSVRZWM65aP5ionvbOYO1WwNP+9FdFHrzqpxw2j/kBLCjLIDO+jAczA0q00EtlIc2rDU0fZi4Qwa
Iz9tWSU3OjXT4komsIcR7Ots4waNHXGPE/wPinzUcSMJCp1sh/y+3d1cqdOeQTj/kXTXU+/SfCjQ
K/Mf+7VdRTVYGLEgvJMNBM7IXPkrFshrgCg4QlDvgb4Yw6KSI+3SXRv+zVFKhJZsjCmjsIBrRt2U
NZKLS1El+tKZpDPFHVmqewrFocHrzi4AEfQZTWYnxgtYme6gXIDlTNqdAFfYUcmPmo4zKG6LQx6K
sy+IdX+03HvrKjJCcaIP8FqefBS25c2sral7kZ2OQb6TX7YHlKfs16mdJWBz/Ino5Y6AE2CjvVXg
t+R8DlDBf926Tq70S5rf5RrwfkIkzd2SOSoA2mqrxDJVe6yzIZ4Ktb6n6Y/i3M2mleF+iQbVED76
HNF7by7buuDl1ZcdWeX1O2+tizJbTMB691oAGG9BX3wvdrpVzOx1b6TtQU7DrXnzxdi73ww9hSZx
vrJt1xO8JEZAxOmlrpTOoqnKr7Gwn9olPLUS4L1xfnl+ACsaIvDI/klvVLyHTB+DXaQc8ywPR8GF
q4D2RtvaH98H50F30XEBZUT+UyDx3zL3sdO7hKoEMF3LsxL5V6ID1qOH9swg7aRcKe7AAAbQB9Rg
gPMpudxFJi3ma1YIqgBNDNKyZhNQs2rLwrw4GH8OAP5QfeypkHdu0vSxm9Jl6iNEIPNLmm2oWshY
PvSa9DCjqEa5e3X5YIIlwq9VOscGGVlUAzRvkNjnd0Y9kLNRpR3gqWhlGmqbr9MV7mnxVH/pfgrE
TfybXl0AaRCLzASrFvJcd8gv26oIAqA+HSJVJAKENNBXQOqROnpHx9ZfmzzPogpuNdfGr3709VQh
kJZ/5Os5aKeyI1FyB5hB36stwh3CQNuZ0Hu+KLnfwPCo3iq3SPnC53Lhj5KZ5UEbgH9S8V0CsSae
L6HbY+39dXvf6o+DqqF+F2jjzX7AF87u8KHh4TMPXC8M22gTdC0hk3mVwjf3/aoJMUVw+V3Sisp0
QpuQKYFfTMNYB13HxtduREYanAO7KQTeYOJD81ZGAMc0ymdCkQtIfDB/P+kY5dP95nc9kjT1aUNd
htDmhyq6GmQYtElfpx+uNW+w5TA2A9UoFAqn0FdJayHv+OqiomYMkfJpN+4ogpm4tIWVMyzJMkKG
FPyl6WmKJbJx8M5ZpKMGKceTT62222NadfAcaiR+NKHapSHrjBOswy6BpMS9LnpKPCEDLI9p9inl
8P2G49UIQAlDXH0D1nF/L7qL24XCWu37PvRMfou+0z3T0lZ8diZpcvdcgpCL+hyGEay0vbb6OBI8
H2gAPrmyd98Hu82khzwK8O32ploT0oMUX9QLAWu+20qX/qe+/h7Y0DWEUtJZNG2GHm9W2S8FVIx0
jyJ2xo28bbTjZ1bmQ6028kdsSVt1sXscj1++YollQv7WNXE59tR/GV9nj793B+EwMooLG7M6YSNq
qY7DKm7SBHS47t1Ite8t6Obqp5eNj+9NbYNCdVWCEHC4Cu2g5NKdjNquNLQ056KeV01Eqy7xXXzu
luYaFUO19aslopAhoFmR1IxHt0kFQXt+u/ELoTPz3iacL+QH3kQ2P4pWXf10tR4UYb0LfvE0vXLj
phrN8pFH4RASKkhgRKD+NJXyxUQoMf+oHl6wGXjJ60gZLMZBvDH3fu69I6uYti4FN8JMmh2xqaOh
6J5Stti6aUEbcAZLpo134ENj87CJqS9eLamY6naglx4chk/0p1Jb9c+wxWEwjuecf9qkwiJI+0sV
P+PvfDUHr/ukT96V1S/KzaTpOWCrVtRBpOTM0GvQxcz1vRpHpiByqS3C/namqvP5Y6kTF3e9/u8a
dOUr8/qiWoH2F+1iGEPz03Z4X+pB/EEF2e4pyEYHZjWCeenx7nAHWao=
`protect end_protected
