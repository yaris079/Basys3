`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GCaPNEXpfbz9zLjkivxo8Xh/lh+FTFCqzE6+spetr3KusXT85aw5akrbtYRDa2TyyFY3oWiC/pWb
WVp6MnAIPA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Lm1E9QKgo3e9rthKRQbbeUJ+zl8sz1tfnG9z5+JOfGrZ+QLOINTB7W/S7RHHMMAkexmB8sYIplxK
FF27kL2MeS7y4Af179LvLc2T2nu1y/Y3hzzkxnSsczaLugo5iVI2uIlyBKyFgF2b9eiNmaaA6Y1U
HE4hsmn3XuImAwZ+m5E=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PuXNs2rWiVl4KXhZUb6VBoQspytDJQnJdPGI7g2IhasUGKVzvaGTUHzoaAEusOqVAZb1mfXyEum7
1vMsS1Y0m+3zWgQFsWNqcFRfVZwdp4945fRYFdtZKDO1hSBdCwHPwsLaH88/UmKcfZ/5VtgQ/3lF
xV6SpU1pBKVenEmDs0v/svBYrc+zwAzLbuq4nmnhSJkJ1QBFk2nq48GRd5VNs/yWo5MKnhZKVc5M
NMHmskEZtRyWTsqI/1VFnGKSE8L0eDZN2Y3z+647xd9MnI4uus3oXE9tQ++zZrNe0+WrmNX8zVbu
TaFcI+HpnpM9uS1MAF3PIW0OBxL9VIWh9HuVfQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ujb1iI69lxSWhRUyEKEsvs4JtLawcZ1bV/YGzwyjFVJy/Owbqo6VoGPnBIIzmQgdSNlQBFlEFGTE
1ulctWfmRnfrIKlPPEr3pk6r+mIWBRKedG/ZUIZVbMsH3Ls1TSxGfCKfHiKtq/QbCfeV9EbHul0o
+f3erXcgAM52mc3xwAI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A8465lc05SLu3FhsojgmKBB4d4h2UCn08rF2dEx3ECHbt4LQRX74qpiujQaVrIcgXEX8AxDQjC31
neYpSrX78k0Q0ge58AryY19YEUV3h5usx6usbe9/ll5UabMLCdQJwVlrTEWQZaEuMZv6EKLLOT7F
6FeIYU9xVW2C+XGFwIZqZZog2Lox3sHjofWTSm2vu0EOZ88pUy3kdQMrZGVfhOrzRMtu80gC6aNr
+EpsC04vLsBLHxSoCjiiYiRtLfSommw5vfSUCvJ6EDvF9G2jZ70GB+oiAFD6DQLStBw/5Xu2q7KA
yLgPxc7rc+Ga4aNU9C7I21a9yzo6xomazX0Ktw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 18848)
`protect data_block
ljP1FUzMkA/g14wAKjNorjJxIcYqvxA6/piL4kHFNvhiXez2o7h12onpTcNmbt5r+0PELFIB5b3V
0HPV+ebzmWketll5rv4zYUpx5nEBclMh+2iMJFl/SjT45lrPuCKrFZIJVOAQw75qHAB/WOtNRbIf
gS5L5w8LmTRd1HPt8ot3nRl/9ixRJDHpCbTaChtjvAUlB3qF1lQXQuzZA1m7mzYu8p1r82AUWW97
jbGVku1sIc4M/OEcGmVKgSFV66jl/ALGUobSy2X5pLeuTB/ELLfKLvqLIbe3+n4eRWZaw7zbRMHQ
/td0P9OGr6DA1uvh09wI7nb0knCuHcV8LKOpLHX5ad9Z5NQIq6m3MB8WRkY7JZKJzJ+6b3ZrNNye
1Ech1CpL/FGDLKCA7QSdEMkdWHOLM15naHMb9pqGTI91vnnSwKdB4T28AbL4+g8i6YAlwybL4bOe
YBDeOPJKXxYnnVkI0K8cbbEK1R8/JBbgA3LwYdx2zkm3qhlGVPJ6+2gZnq/ynqiCnEoyhJdH0nLV
sXVbNIjxCHtEq4fk03lo8meqkMvnY5ZeqeKe6IwbSMgQizTra9B74d2cHZNN8oLp2lG0EjNcRHGj
mAmYi0tOlD0c62FIOFvhm+/EaB4OTQ44j15lPq2Akuq6E7mj6J1vuYBO5ET+BToe1Mz2hFqd5KG7
p1Otjdk/wLQbF+nN2pXSCMubReyQSSoeoNIZPtIrt8sL2IfGpGsf29SfhM9JexT7gGIfxWKqIX8R
qO+hnFYC+rKl9bwAgsQg5Gjt9p9u8xrp+VcglYfXsu4iVIfw+h8fc6pfJvwBIZbFSSo70r7ZMic3
0efp2pQ5G7DZSpot+JCy1++6SKLnsnJSqrT54VLYmz3oRn7JLjO5JWdXSb9Sx3rFlUsXNPsHjvq5
F0b9n4uq67a31XFhyTOlAbrJl8fs8tHnC2/1JLvgP/mx4LdaNxy2PFHlS9OqyBD719K65s/ep2kn
JJeE3giyZK39q6GDkjpjKflwsgRKjOx6/VCcNH4Vbl1umVAsF6JGdSPvEwjtWgR3t0EppdbxUPqE
aqat4dj77hpfUJ9STExnejtv2r9CSQhnRuM2U/Ut7EMjqZt/Z62IuGSrHENeEUAmpbRWnBiNgAao
PHOlPpZtF8ZIWcHA0fAj3s6nKnWewV3sAbNG0oopJeRlTXXJTM7QLl125Hdod+kQiITkJOzDWYcU
rlwnQOP9GM7J1hsZ7RkdPS9XSZRmnDnK6JCEHV2ScK3WTwUKcUpdc87+4m3TdAM3FD1Rzi2aWFVE
YlGVZzzNfdvcxhzYtucs98WlwMs9FkmFqYSdwOVoOploCPxTyeyCTvX3+xm22g3neIY+T75UZA7T
Uxu3ZUe2UC+rlIz8hAiPIIn/T1hmfnEQSjEa/qwvsCCd6DyKwDSTaJO3oh7iEbPswAEzUz6nOjTB
Wd1e8rBzRmXr08maLjUbYQdtr3FjD7yDBGPkbJQUL68JRfRo6G2dZc7sDyBvx0XW/X0CNLIdrmiq
sUBvl/OWWkQ0MSWsoxgJPoKVg0LA4rV26qAopqXPDQinW6q952fuGONjrjwAP/BN/zwTJ5TupTM+
Is8PkteZFteo0cqLsi1wcR3T+PgE95HJg2kB+KZ7BMTV2GhSES83sznj1F7IHbyw6gXDl9EdgvOt
K5aM3JZMAIrq4WjZmHpYkr8GLJT5WIidX2WOeaacB0qGGEIHI7LpFHFxuzMLs+X3svgS0/Jm6yFl
GKY2fdp6Q7xTWEe8atUq7UAgLRt+UrPjKDBZwG+rD++gyu/5RMnN8ceXOrUJLVWx/0psPG9oQvgI
EgYbze+Xfu9xnBodvVlp/9M/WCYCg42DAP1ll1bNhh9LkmPyDTnCmEcc84/A7lkFqMVv6+DHz1G6
pxC64MGvFl4ok7VnMffOaBr4c+UMVtdXKlWSeRIlD8jVyZ+AYjQssXXbQ1TvmPLgjU8izUzHX3wU
y7weAR6ay5e640pn5KGMT1KJ2kvJpInN7yT4+80YQpDp+0osI2R+k5p6KyY+edwAQLVZ0M9e0YzO
FNR/ZSdbhz4YiccXfD7pSenovo5IUld1lfQVTS/2ustZzc9dkpmY6L0ziD8xYwItx8lia8A2Ozws
C8UTzzDT9D1h1zLa9dZR4LI0bhP/DRrbFSgYmUJqj52WlY8Cy0zxfLAoGW+tjYKevfv45f4k+/nt
9u5H6CMD2kJ/tif39+jF0x0a4Q15IsFeLArPjDhsmCm5sIx3hY8fPY3GNPxiXB2ydMq25br0kUXf
62HxNdEU7lZRdOKp1zMLr3Es37+jdh3J1DI4/z2s6tgxv+Y1VbHZfgRxHROyOc2Ov5fS/lXCg//t
NyeUiUEmjCdC9ERE/ijsKvBCqdcvHYtcgcAHsUC8E16kiPNGiHOAZ/hoZZ4nXEvpk+pNU6+oQe+j
VQcw94nPMZ1x398EwPCpbM04zUcIJ/ymg0loUDJb2ll0h7rBc2o3RZ764DjsJUTnyfMZPdNbOLrE
Y/Z0KPcKnlFoBPnBeEEFGvYH5GCzx5z+MsJ6Pk/DiQOdIvj6tR8j8oBSbGVRI1q++9enkQI7D8i/
BslzslaQmEegR+yY+ourkEE9BolkF+GFDnW3iPtqxyjNxksiDkQQGpMSKkY3ajrwTTmdb2LmwOov
AzrRYAmCYu0QdCJ7+hUbdAPIK9cMQPv+xADISLLpRn2YggMdX0cwsseNS7bakkNAKHzXPCSntNTR
frj3gjnBqFMy32Qb3EKdqYYK4p1r/ra/nhb0xJT0j4nQgLkB8rVpenTSuReHMT7mvPC/T7miDnHZ
0xEONSDn8xQ2t3AswmQgzTWoEnhf2GyPOTWWXyWtT1a1M0WRdqDDWNWcmU4FhxZl8Z6TvZFgsKJT
eDrnsQE++WnKAmj84bolhNc7AMKK0o7XieVAQjw4802H5NzRcgQIaQ6BgTw19RHFiGOh/AtfiiIO
Wads2p1dhM/xs0sYJMRDoYAy5lhKeMZjpjcQGhKnrIerWRwriluUL4yfF3cMUrcyc7i3c/WhJJkx
DogtUvZuNanQFnnxg1GxGcH5Rfx3K7fMTBjxF9jvCPcfZdQ9hgLipF/s9iSqZw5c6eDABJio3p2U
qPnB8LzfkIJDlpTneqblOTWWtynYxjQyjaELgDxBwOTJjB/nw502i6Nxf84OCWqFw/4p1cdtPxqQ
tRfmYWgfPA3bKRJvL9pNsEx2tyNprlyI+1Xe/GTn6iL0ryuWkFQH1Vn+DJ49na7kKlCkNQovwmp2
lsBuabTEKi7bEk0mDbxdASXCdaruvb8748sRM8hz5K0xfOanLAj35Pd9qyD16mRxzcT+SNG5jKfy
zocDBxFQ8zmxKNfaFWpDEbhTvwX4Gpb/Z40Zhpnk9qQLV6easdhhIfEvd28ZIruUpLdB8+j6IS/G
VbZCqydoZwELLd8HAhkYKuRYgr4+JB2qvHES9Z7OWGMib+P58OZ6+EabpTXAfoWcCIbPzVwPtf3F
dy8gJSbwly1aW2cgSPih8xi5+WRryuGlSZPJPYxxTHtvgHUWztC+TIQxQnHtfGEKp/OVuLwV9PIq
eenDrgzLCuY1x3sKJ88vj+gqoKx1w4YjWu1Z3TD0/U8S+8W4HscXW23jv84lTcM43Fz9Ie0nuV40
dvn6NXFui9A5AMld/qKcFHzUR9AdoCtsT79P8U2Zy3HAyrKZrpZAYIt2T+MlcyJNfRwBGXeR+U3s
qhLTy+F1qPivP2dXF33wq0NLLQnAVFYjahqOluHiFksSDFCGXfJnigsI692AqV8OSg8x2VEs+28p
CFkzMvtXAapOqJ7czqk7RzKQUL3Nt8RgTa9SCrvLrbLNMWjIXAhAz+pYEiGWN9vOQ7Z7Jw8vAaP4
lwpbkepmC1v5+R8RL3FDFdOpQbCpleE83vR4eXFN2HJq3DHm+Wad1G7/JGrpEwwt4umJFionveWe
w/Pzgev/6IYx4TpQM3W9WofFurpQQqRuMxQ8UMPgudELvWyfFnN4HTgQ0KJibGdsFAsCLrrp6Hu9
yfX4njJFAL3lL+mDdRznzeds8kWpx3UDFV1MdQWAFdJr3z5HFwYqu9QNtkmlVNea38uiOQ3fDtVr
cI0E/DO9smQ4KkfDRwFery3xV3nZWxX+DDcNxLkBBiHCpnFGucyDgAp2V81yrA/BBO7tbV/HjQPz
A5Ytm+OvAibMO7nJqzZZuBUSvUtifuC7MWpgfPvcSMvZxyqz83kABrHpsgJUZNDHN8aekgMiMd29
/CM+xcTt9c6ELWZy6DRr7paQbImBU+AhjTG7ScQmipgPteCfZRqdvstA3NzwvsPXwsacncEWXfFP
1eTiy/NDbyBWIgCW0zCIlVC4up4UDG0aS7BCbHjzYz5m0bhqFvwvcNrEWEaCPVRha+lmPxkzliMg
80cM1EtnM6YxVPkLULR6lZc7i7JjzjhLAx6xrAW1P+1sW3X8APlOcoqUxvCg7JvpGnkdtrYF9F6G
D6cXgmGpTPHCGa3uUo6ji1qdG8wsV0yXAfKVfjHNbryVz0J+vDK+1kXPuZ61pHljqwWZIKXQMe8c
7HN1/Mw+WQ80vOyONh4KrSb97gQTwFzcoVKCz/pEl049QT101FDsxC0+ZdwhFLY+ffI+HIjAZ7wb
Tms+1JeBKEj23VWTJqgsnYKMv1a80CWgB/bCBZeFDSQ/CDatXt1BYN5i0KJNH9rvnkBlE3WGhraj
nj9E5kGTgEuRQKkEkUJMj9Dje7md/3AdMw/GNkQYTUBB90F7cNssURuE5AHn1wicy8Ul+nYZChnV
V5zxD3yL4ZCxUhmDIzlz5LAEFm/V/2cAhSQazIwdBhmepnA0pXsV9Dgghcs9vI15jDI/Hfc/yo2T
LojscIQURjzKgxpAgNklrBs8tI5paH6fG63IgUE+aWCq+Q/I+CPjaoiNou1+7cxUMfVUS0/4Iy5h
ndf/gvzekWt0o4DAbzNX/w+nPoeVd5qqOAwqfT/YbZgghNfEtNVLpz4qmX3Vf5gGWYaHnkG5MOdr
pmVZkie+5tXog5039tjT90+bm0t8uelyd5E2lkzgPU/1hNjC+/4gK1IKF1I3+wO/rUHkhSmS7fVU
99nKJCBiRuTAsDNtbVbeBhMSqpDZz0eQi6pDq7z3mxFCUzdIuO3Tx9e8466wjAA3rf5EcG1FzizJ
uKPyZjOJzSCE4qK3sLUhzGIj55VKTZgj9WdeBUkxOa8UnS7qZ8z5QizOaaYUzK3MbGyP8id7wm3z
gK0jKQP+PmbTmMW1ZbdU/vqwszN2A+2gAfkQkDUHpsqGh/IKmO6QGLRv+pZKt7q0jWIctQrd/CkE
bgQE4WvmXfPvgpzAAmnE/UYxbFjaBvTAk4E/EwLxA/WBcslTMb9SbHrI3lYbQlL/LmlWtUKsoPuv
1pOQIB8ObYABaiNUrswPMlXZ7HCx+RF1HUNGiVlcVxo+r4Sh0FDzyjccjVMMc9LyDfV1JFRcZdxR
1GJ+pD9FfaYigB4K2iziIa38ShDrp1BljzZyFebJnTtDstxkB2CtHplzKTQsmIIomzniF3mr68hk
sKpdu5BgY4rsGemedZZ8TRWbW9VcT9k7exftNk37AgkTmdiVClBGaVFyD0kyvLsmU0px0Nt+rFTc
U19rnrQ93F557NDwqeJ/OlyG1N/BqDY9ARN6wtXOWozhgsJGhbu/e3K5A8BwjXcs+IzKlDs6hV+C
S+goG4LRVK/lCiXEmiIq2B4o3yOal1/o9wZEOg3SogIXZsNb/UGe22RGdCN7ZOXxU0DPjpLt/IXn
f4AhApjtULwnmmfBez7aPqyYN3n/LlYBXlS3ofHUSYxxKNbb/oHFVnAgM6rrvyvYbT08jJN/sQdM
NC0LDx+dBNoBsteWODD+QfqA/Ua72nj63DPov10n3FMy2QaiBcP4BnbEZ2fspiPqAwkIsWDVfbPh
5U1pI4h6RVP41op10Q8Um7PB7x8ZFuMMOafAwnw7SHKzpiSvojKsMr/X69jPRKyJysJcur9iqT6j
2a2TyCDy2oB48HAru4NwFmydu8GG4MosrQPLiulAiVZPtYHsm/eE/1Jtkc/gzV3xFwOb8KZpPQuE
0BPP/rbvjLgN9D8InI39HhaoHc/quR9Zh/kX1ncJS+ukdDnxEMIQrU0pjC+60b2W2U8rAnNfUD7O
JLjYPmxtM7IpsB9UvmRlnpBq5E56QXK3k8LX7oFQRGT4LhNYqX20ekBd2sPoun9eoozGyC30iW0l
9mknLgKgE856pBgSWKGHYtXYjw7I3a59s0Fr/OSkKAkvLEpM5QnA/wt9sNGN6rWY4akTX6lK21uM
gOnUmybO1MJU48/XgdsacxAa/q5HflcJM4c/lnN0byjH/+rNwOoUn5ZfQtvAgtDd8p6cocXiUbc2
9i2jBJCn0OqDPYdYY+LJICYwAaUmP3Vovqlc3678CCyCJlE3kcLsMxvI8H4wkjsH21/2WrRcifEL
P2nXGQADHgG/6hTuJmwqMPwDqJ7VimZHacayRNy6UZw4Lg6d57QhLOVdGl/N4x3wgB5UBHUDMDVy
7i67RiORVO2cTJLuhzIl0JqxQ+2mAhkDn1KaXf2fDgxcp5thkUVNtobZpw2ugKfLL8PapVpU5ke4
pUMlH3E7hPMz286Vrz/UWLCPy6vefYhFtO8eFhLXnwCK05/mFIpRC6WVMNbpkxXSGYVNSlNLpl2e
AgmWW+0kNF/SovOUoWsL2r8nx6B0yRCyQsabZfbbpNIw963k4NYsUMatKWShdRn8aU8/M1B22BeD
b5M62PgQ6l/FvPlX/AVgmD2i/TiujdHZSTl2OxxDIXHENE2cQrlP711wLW+9nhn0fhcl+HbVjhrF
HVt9emYhK/14UX453i0gasvkkhcHmhMZpIyFWuWKrvXQs/348y37CNgwSFcuXCYBFI82RnCJ6w/F
CDvbKG4H7c9A5RJC+SoV2BXCak980HGskLnj0IghIui2Gt6HsqFluTcYDwo+zy5/rD2vZGJsc6G8
25yamDtXhoE+Z9jHwhlGfhd+pt4uCmoA8rOVS8Q+n/KEfbxquXa0TS0hRZNeZ7zAyj9NeuM0cxsu
3A3IeeW6dN2UmMZ90KCpSjxo27jEsxMM7ifjVtEsEsy3aaTujxExOutl65gMKrJmBREpN6/Rn2QD
6pKhzfK0o6LpEVNBx9NCl1YkLbbA8uDt2o+lqx95E2DBStzcQjtj47lvuUUjwdtrR0zmgq1LHQoa
V7O6yGjpfHNs2/ni2am3m7DJQlQJwTI12YeIOjYoUSuBoAJ27tzN/FU5TFF3zHW6ffMcIXkKzuc9
lBxZMUjzJYuLPti3+ZiUhOCxBRCtz/AwueVW7B5NnH89WvWzfSTBkLptM9DAMVEiu6lxBRAFivLV
u5gw0zYJTPscRZPYWbBmsimkDe8/21i64XQaAENkuk+2qr+Owc6Fcujk6GqSegToOz7IW6t4ddus
fizhkecwghJkCw/HTZTy1luo9ToeLG50sZMRC9loJ3+Ib9Nn3BQuHoemiD2W3lMpoPPAsMC7j2TZ
e5ELWtbU1RtQhTPBLd2MbjNtsA4ObM3QkH9DAmunVXdRiwWkAkrvQw17xDmwPmkZEDRG3QCBs8Ki
dCz4XoJ4C2mPXi7quiXx70i3jxux3Qz6YcU2lckPWdvjkrFyW94JmEUqvgkcQLkB0ef9k8w9tUUJ
7vzXBZekcy66OVstN0SzUkchR6Ej4B7XuVtwm85YTax4TXEJlOqib7FKY2+Gxyer25w2IYYGOrxO
LZLpAUTsmYlonI9ur7sLsSsNthO2I8AIqpmRTzA/6bWTgstFt/B1ZLX2GUAKUl1fVTd8oIhQPzLG
AXMZLmj7SQDszQ+5bfwq6lWkRGVHq8juIB6xnHAWjmVVRfX6UbmbBVUIUL+7BVKJWa27c0xlDVdD
vpj2bK9pQ/VQX4cdSlumJZcZL0ojrE9fglclCrRFnHg0XNUe5jvAl2cfazalqbusfkw++dvUEk5z
KwuQRb+NC4CxKmechwZn8sA1WqU6yQCPrnbjlgugFE26nquLTcTfxw6gqV1F/NAvQ98hAe4CQchJ
si2v6nteSoGBJJwr/qcBTs77YcmmOOv9sEuHnBkDHNSp759PuCOOnx2V+SXKORIEZEtSGgoaScRS
bZIZNMYSMjvFNczMMcc/eQ5RzpsGvmhgEtyFksm2saS6mn7R1qVDJSSYgTU7u/4S6u6u1aH2B0em
C3JGBlaPWJzvx9XRdB/IVNCfh6TySQWhXdq/tua4XQo1MG0032dTBgattNyx9rabhe6KRKyWX1y6
+E0BngZbv6plAKppcNq2tEJraQv5WYagf/at/SzMgUUTIZe78kTnBRLWWmZ7AW84BGcRcciKzCKc
bHDgY1cPomf75ZGdubk+9QXHGcRY1Q8lNJP9wz8B7NNg52BSzEuncXTK43p8EDlLBzTsp5dIcS10
OtYxOO3bBA1o9UptS9gO1V7HSNIr9JcvCRR73Om0Lo4xz8HJ2lypF2ukjxSkMVXYXNfuUF7d0rnC
bTaL/wv0NFQ1WgljzdNIMNi1q9Ti8BR8fN38W2KJlZLQDhn1YrIFGtzxMEU7vOykV7g193qSO/s0
LZi5Ff8XrD7oE/NTMrQCF5sQxaLkK4O/RIwVw47YkYxdQrD1VRuyqfYu+DoNv+mMyi/JuQdSFRk9
I3fSJq4TsqG4Wa+YaN1iRQA7oyZgBbm6yZY3dcuhE6GQPK7skxs1pJJbX4HNR+/hVIpX2Txf1Iz8
0oIuS8zkxy5RVF4RKQ0LpEQCnVJkbE2N4HJ3v7b59oaX4fsWZ5yQRpCmTzybwnB8RI/Bn533Sopa
rvErbM0T5UwBwmYo7Q1cCaLYk4DK0AN898TAKBejxIXrA4mreXiYomlFJAmicNkz0oCpCTPu2Ysm
f/fdMK3YBZyyGp7mnymWPkeTjd0akDL8XfE6UdE04n4NiyixdaaYfoJ/b7t4UVnupM/AxY8yjy2j
yj31BW8QgIRI5vogRymfkQJ83zjbr3aJ3gZ3aSCabE92hFRv8Ly+pVwFbr0s47eZ3zgZ9MxFOssz
8di+6Nn3Co98Xfr0FJNedFSWjj8IjEBo3ysaUPAB8gqsAp7vgh9Sci3KsRk3q8U7ziquwYSgZ7LD
OYppcFyhznSliryA4OAC9aQ2Zbl4ehE/8NaVGMIWmaN0tHjhKIS1sePjxKNWPDGAfRuJ19PtAFzq
XE0mcUet7+ETGdRQvpYQHAesBWgTZ9r1PW1zc0EQUiXfM0FET7OP35neO8Wj6AMw45W2exULc+va
dbuRHc5gZMMc+1KvqfizkJuDcKKCO9eosnYxJkPPFgTIKD1yxBi+QYG6BMVnrfJUKqrLANhsPTnv
sBXFyEkX2D0/kRqWmhpGC2/zETNx1zFL1aGPdONjwYWrcQB8cgCHu1i3xCdwf4dwbAojuiVa8GCE
WjwloOWRwLQ0MIxvItlA5UDnCuDIOviqJ4VwQrDIYlpNM6cYiBnHHjUjJbsznsgArTHcWLd3hfUA
tUpGfe0c8sWx9ln30b/kCKBgCgZjshOB/51fI4rsfE42a9miIeUobPvVWxpDxuZ5/OTQkAAB85O6
fedeO1Q+M4k4PPom+TzIxq+L8nn9ZWOWMDe8VNDxqFliHie8m6OUFpJTWtufT0f/tQFpkwl0s712
ShyG3ylyGNJRM7RVGB31l6e7pz88ovxWLEdifakTM8LdKkdtxcjSChCsdudOaCx+jL+C6ZQSGhUb
qOgCzFkYqOm3ld4O/ZofJJTgqLPE/dZrfuMcg6wNZPqpcqBLo23nez2HbROO3tjrkV2Z2kW5sZm/
3wq13Z9bcs7G/C9aVF5haM5QteNzIFoqr9bXoCr9i41qRStatnAaIEtanNeHzNxlY3TYrPsTCa5j
YuDKOfflK3Q4aUhoMN2A1Tl5W+n/8drtNRMND97Z24Udu1tmK55Itnq9CPedgjoLHQKbPDR4S2UJ
6xS6ibXE+grn7orte8qEhKdSPm1yRxJJwjsyiL3djVc4lAD8lMk3Z/kPC+TwFhPhZJJ8D3FOBZgA
5I77C5oASdcn07DhhKEcIUoNrMHuzpbXoL563XMs9NJXoWPyXs6sqQVSIZaqoK/jUCXmLGPvPFcG
1CAszLtXGo78oTpfRwH/oLWbGw5OHVbDS2eZntUFKNNHwArqrYk+tmU86Q4KCY3krUdYcWZiiAzq
kaRLB/dJ9QMRUWafpZ97S5ukWcUCTcTYSGTIodeJZt+hA/Zv6fSLAMeLo+iTzogiQRsjT/KsMbTe
I1snMtFQp5pAaihpwS5iYWGmIWwsYmJXlyVE6MBNGeF03YJhDUmh8hbGPZFoxjpIoBgPXFEQTA8v
HNf11E1gw8pDtWbWpiva/kLPRfRuuFKVlBJ4USvorCdSB/NDQxcMNj5cz3ANY9LEoCw3vEloAmJe
fB60ZEv+R+va6Yulrs8fdMGDCbdpU4Ox9yYherH1Y+dvTJ/wCcFaq7dytVhKtXS73XZpdrqK9CUT
V0pvstu0eN4vqgGpR2GDZqNiGtNVSWA2cG9a05bj0NI4KJrKHYQNrm+Yc1TK+HLTRi6nBuADC+ij
gWMqG2zul2scetVQMx3D296s/RQqi1fAxo/Fj0iVVcLtxD/N4e952gyoTQFBJI7YE213dsa35lz7
IKz7pHRyDu3EdIxcQtC5qehPxkxIJRGwhZ7PTtQNEZiX1pEiKSyCMo35VnNl7KRU1TvVxRshv2dA
xub0DPdAXCUTMZwePrgBA2YfN4Snm8AKlRD3HoEq6MU1HNucwaROKLGAX0G5rciWmM68TvlUdnHY
Tyv+LjuZeCfalHaA/xWLlNHi3ZU8SJ6AlNlB6orQ/ckBn2gKnaM/1qsUQEiywO3pYUzctfUZj2v6
xvChSp7iUoxE+HJyCKl0WQFwN34CCr4wl7qMPP9F4EUyUivPEEi5vjisLPkpmyp/h0e6P/k49MhY
Fi/1AEt/ALky81wXEwBxGIj1wQ0ep9ILIRLejP3CTlCauEqpTVja48+UFP3UTUcaq4b+S+OOu4fM
4nRpOIS8MrehF7mKhnN8OK06CsVi3cj7YbchV3s6Bh9hcA4GG3IBIjnb489cJzhwIYE+FgHeEgv5
rE53uGd+jRFh0UhUtU3V5BROgbdGwJWsQz/fTds9tQNJahYc+nhE2YNPY8WUbiThnnjn044yy/Jf
av7MoXEJPR2JasNz+cLKH6C1dauO16AK0HylA+ZTsiUemoY8jbq3tGm7qvODwoaoXw3cKd4fzqAi
moPXG7pr7XD3q8Yr01QaIjQm8l+xSna+P6n/Z/eGyWHTzSDU6qdDCZS1fgu1y1B9WdSYGh0Q01EU
UY4Wdok/pRQvxLuN9NovKA0EQ/fPOz4DnKF/OY98l2Te8ZU/p1M8mzzqivmbgoOtz/dUnppWsJ67
m76fx8bMc9iPudWJnSNewB0m/S5hhhZW0nMAmgegrqNXyt6/SlXKWLBVZSUz2Juxp++7EWvExOdB
y64mmlr/yWF7eKP2Ci0EfSEdTMX2GHDK2/EYsZKdwsWuaPV32Ve7lyVFxflJWtJI66CUrYuQkXb3
SVoPGCqQSwnqjYBtTO19ylKEJjkuKck9TPiyey9fw7sJW/0ffHCYb/D7/u5vVGY20r7ym1iQjaY2
7NDcO9k37nidIMksTu+ELbG/4uZZAzoXH90ck5y1qTgADzx7YIpP0GJwIsZNa9HuUUaaEJxSXdYM
9k4AtcC1/gzaM/ELulGDupGYi8S3fA8CoxVQF0GpV9o0mRHium9sharhqvUTMQCxE93C0POXPqmD
YcAf/9xSgrSFG5lo2MzJKOO3LJyIIuSFAW35HzoS3vGNy8ftelLWWjWeZoOj45FqzPFqFBFhO4vG
RkG8fosmrwyuWQNHIJARgYQp/0prJqkc5v2peajB07G7WdQMwN8P6NFLaIhBuh+iq6RewHEuu9pP
1VNazH5RJijiuvAKCNRD6g09Ku54eEvEqnu3zduLI8ig/xsT3o8co/Og55sum7dOvRzDICHYOsjQ
gwFrGYrCo7mNSJ7L13qTKEt8AVk3LPeoDlOA7tBt51y18YeS1Sbcp5UfIjz+Y98Xnt8RWET4ch01
HlAoO+CaI7Rfz7C1Crmzeegv3bUu38RehChbceYuZPCaZq9PtKJq2OeJNZ2A9DJjHVw/0PWrP1wW
pK2JCNnQzyqB2Av6G2CUtvpZUK7fW0ouN0ZAT2bYoGnEry01mQyos9WcDrazlvTdZ2uhNpDZjOgt
WtPfmGxHIDeKEBq973V8HFDVGsX8cxc3fDXdUjfSkSooOUnJAff9EKCD1v+WfzSbemoI1uiSFFYi
iG4tAUCp3VUreThMK0eZxUjNqeubZ9hvDOVV/1O7rOlUdUBXXq7MkmyRuyvv8h0KQbAFhMR3HaSF
MWAv+P99t/rH8elqOM9e0jv0efk2Ohurovs7IpHeZ9QwSX9MmY9c/gG8Wtjp4iG6cgL+lcv+yfXi
EJrzMuvYAB4Op8rXFJ7eCtTPWEo+Iso7vXFPl3dSv5Z9Fcb4BFntGcGR8L6dGIrkdcxrizqUDukc
9IWGnSrbXCytqIPUM8uRzh14bqeHGb3JyCXoIK1dXzEP44OS7NLoDppNwm5Nd41YYCvzYntCRi+N
gvsR7y1XIeZU7vE940LkrMf2FF/ToBZoRag5cWQIbIgcqk+/F1gZHkkQFjaIHntB8/LYQlgDQfac
pBCZs/wgExynhyqfM7qUH5FqvtYRa0RE563t/XfX/np67xpIN2VOXniKYAQblXVX0Hk8zoEOFWQ3
VrRh9CB1JyeAWbzjBE6mnU8MeI9EaW/5ppmz/M95VFraQ0jeLcSKoj25KekDOeRx+zl23PhIvVWj
xzQ7UooE3HrP1zE4qkJgYmY5jJqZugpKXRvfgNctOl3/L0X1U1y38BALk/clEM4THRdoY2mzftnA
R9cYu93oP080jSuEXJMOtI2Fs2nWPDTM9QhBrb/EVdOn4jFk68WOmKM4NR6HwvTtNyPSg10kmgcJ
5G9Affmzzr+6qFLy62SZWVG9BPGjkl07SGcbPOhjKn1A63NBzUuVs9VbLaBGzbm2xnJ2+nMs+Qyd
w4XCo+M/OonNOQXPcqW9d+1akS+YsWNNF9qJvaqvCc1wLqZTrEw8nZlSl5v17A4bcab4OSA3ZOEj
RWj1490Hj9PnoxoraV7Q/afnIQEYtKs7EQ/NBl+IYOkRvmcqkJQ78sSnMVLhXJcn4uyvoJx6KhER
FS2jwe1MLd0IT1wC68/mI6HW7BVMNYpjPZ7hKXm7fZzwBOAVpNMrjUboAvI7SKRYRXAnAjzDAKvr
jfMDVh4gncgSr1kJh8KFkwzRyzKuMoBv17soFZc7Gboa+PnL+lLO4riBZhCkhoBjVMI7LltodXIp
Uv3O4N2kwNQUHIIl105ymdd7GbM4SgFKHb4yQSLqHKQsxgsEm5AT26y/Fk4R9p3OadHLC5YGs0hC
je59JvWpIl3P9pfZpqZVIo/2lHM6on5KGeMYreSLOBnJ3NvdGYweHcDngjJE8/nnBfTRmbKstc9H
dARIAco7uKcGP6IrwZFSdFFBY0ArK7+G8r4hgZbfZmkCmo2VHVTKndr2ADSJ6GwSsii4XpIZHgZJ
9xqxu7vO2ICCrXAZujv7UrEDY/674sbIbt599yYNHRNzWCkh2G3eenu+rhG0FMDKP2NWfr15pSQ3
pIryPvC/fvNrFEEwFqvEMfNQrHGrvsNt8wML3Z1aeySScDF8EFzzgqRTUXcqYvvYtawiT1J2iOCp
jXejG5UQqIOQSHSUGgD3Qrh9RAT6fVmq9Ovdt8Y1qJq4iovjDIvkUQJhRSgLC7jjo2k387+Imo4q
eXXGqGunR4qhUerAGa9uNIIL7Y2ypAhq4iOXaez429fidG6FTL08dhtqtNNDPTAhkPRMGe/SMRTK
wKz4fLzqOcAr7Dhsr12NBb05XmqUu0E+2W132Ws1cg/UHIr4+tsaEfBZFTaX/4+NSjLS5vG5uGlR
rsUz5smrGtn9C45tkv4px46iwNJtxj8bYiDCGAOmGSSawfBsG7NpyNDtr8Q97RJUJlyoS2RyDVWI
4OxJCTje3ulGUpMITCgFuR4alZd5vdW2KXgUWKibflg6BEiahFOXqGK9koA+GHGt/NuscDEDeuRA
Hh1rkMT+i7fOkAverBg3FOFgjWKiYj/PNaLb5DHqWVWywWo6DwtjCbOtl5PZV0PaUrwOvjtnPgAH
fwW7jno8PVK7OfsDOBS7hodAWe03xJfvvE/mIMT17d25gJliW/9F5qv1oA6nG2HJChlSwmVbeHty
DEN3ZGhFekc9y95AiLeo7ORfNbDX8GBs3PHAQhX85cd8dCISCWnk1ZZtJ7+lvIKxTL0SKw5+QLim
WDbZyE3WC5HtfF3eKRNPl3dGnoBRtvL3dcz0wEy7AHT5htK1Sbr1vkfRQD4YpEdDJTN67pmRhB9e
VhqCXOREBSZhuMsQoQo0bRZpbL4Ct9XqgXXzC9Auj3nzIJYtMLIaqvOejVSb0ABJFxmCvaPmKe4N
5psbHSZn4KOpxJnXAW0lcnF3ayqiJBVYdSLiwHxOkzbvL//V+TP/H2hvgXHLvvqmT4Q5xRezQ0Gz
ebR9B7mNDV6VHazE+qt9cEE0AeAZ3fAe8bBLdeLFNkrj63CAWt0xtpldOg/OPJ6iqpgHskzNzCB1
59Wb3QiTY4SmDVyZTu5+hliz23khKGxD7ryYB+Kw8J7p20O3SbjQ+aFVSzx+mQC1j6aiFj1Iu1Vr
2mfkE0abzf6YMJi/at7cZ0AHeonB/yQs8UaU8IeopaBbh8KTZ+Na3j2n1ckzQ9+aQWdFyfd4Q4gH
CmETsh0FPOY343F469/jqwq4ChwdcgdmgNo/IWx1Vncys/VFqpV5jSo0fA13OLosusKHyoN03Kee
Ock9KdRPJkHJt8C/GeYgdumRM5NuV0B//PpITw5VYh00a0a7hfgNV7Dw4ot5vdFhXr22szWA2V+f
t6hrrmGV+KHtdRto6J/nDArc8QuHgvvlfuH1I0DCUaBdimQ048NooyRDIwoJjG4Vi3JzffYaKY6P
+eMkhHYUy2lcB4SGdEQK4754Jr6S/ZWVn+H32z9p5bdbSVN5MZn83Jiiudr6RQhnoEEWuPKBzfPT
SZBxhzOnBaUmmLd4lqu0YpyNTHECjpfMKqzTlqju5Jb7Pj+2JuXIrN2Wb1eOZTVAelmOvpKyQKq9
BMPFeajv2UbV+4c03D35tjqa5Y4CZtKUPfl96+4i3x8oNA/qSEtXXD4k7JEZ1GGK5DmSGca30erW
/Cpg/ZiPu+/ZbL15sEoSnvoQECItVFenXWySS7hZlAc/sR9SANeSh0odQYXCRst1qx2R1kTCYy4C
IjAI+K/Dn/7V5REM67eVfSoECJ3KGTvwMpDvJNduOJsa0T8d1wbHmAAaWjK8ySuNJ/blxEoZW66B
0XlAwgF2OqXVK6+Xgi0Cs7GI0bQ9hio2GcQi2pVUB97tArjhbjhDoaUBLtfrVp4f+lZONZ1AY/B9
CjGnULUflzT+JI2iyqjS20aJHlo1DZepGCPD2g+KD+WbdYaF146fhMO3B+w01r3MQqIOdyKoGzPV
ulo7qhhNSEn1vSlqPQW0LsA3GuI1fTirP2qin9S8mPmNp6D/ANkIcQmp6ApLBUYTt3hCRUOAWKt7
Affart8BKbMNxBJQnYkQD5ygi2l7iiMtkmvNYJ38BzxbGnAaxAC9t0cVIs5p6yhxnz+8psWmJzuw
rxmQjR+aJGtzb8tRivgt5rbKnJEJ2oFO12pc924GDtB1+ZIyNXH1TgpfR2o2a+Vjb5NU/xKq1XuQ
Sj2DG2ysI3EREwfe620PXBvtoFpAqxQOfI3pIOwgE01OEEMUgDq4TFaY6wL/rj7zLfMXYeVV6pdD
tmKgXwPgpFinbTeuxJm9r/wyJb8gMS52a2JJyXdJTHw2iSFY42ne4rfxKzoxITd0lPWyBWeaUlSl
Yb8BLK+HTAZgtuAi/MpvwCIlzeenk40GJDQ+gLWU5H9wFokG1o2qxtHluYhQ4T4Gicuupi1pw7jK
R06czg8trJuXtlD2+bhm3ybqzxrFLbaj3j1YVOHR5dtSaPWdwhbmJltCrnXPtHPA/LaTcBs0WdoX
LZt6h1YZYS1EjNV5AAxL1iCZplTN26Xqfs/zpF/8JfnmuYcTzsouiPEc0tOpNhzcsJ8IHcqvdh3u
mtBLuMArBoEBZ890/wwuTjDvzhl1q9i9egKUjjtgSy7Sa848DUQFg1AhADeUkc1Hz9ZZkKevOTOv
/IgNe9KQ8wj/iHTAeBiq61y6z0l8qWJtxJG17l3cD9EDeK+qKthOTppP46F6rLqjY8OEY/vDpYo3
8TvPm9DGe+d3oKlCbJeCtFd1eX7uM0I1iOhKWcyKzXih9NRQtBZjfe2SNTatcwrptbx5IiefWjJR
EzbTUQYn8GsHgBhFy3DPGvp6twypdpEBz0oq1y2qkTWoBl/lF95JakhYYnOXyKpkbaUMne97FqML
S1YRolyo5klTY7wPvFhWHdou0RU+2hD/35rtiqC1VGBQpX6J+4TedrlE3JIFrlWlTkkCta6e4ohW
vjX6Uasj4sZ39t8AzjuwTpu6+MO6TkrSILKA912a/FqM0z4Z1AD4ShWCr9CeIHDbmQolNy2otNY3
5t5vHF/wyIgjAOF9qQkWDXgGDWbd8A94iJ/zYplgr0aviPKfg02gsWNamVWd+NFNftjQPbj9kTNx
ErdtX0Gc3truMnVv8qpTw3cM1ukXb6yI7/zVcJtVyo3kGreg9kRjrvBSFbEVwubYahQJ4wY7gzg/
77RYclWWJk38MNaFQ1zgQ7wL3aIN7ddWOvx1UzQkVCk31fytAr+AI1nMbYLxCO4bci1fsJGEUhst
L7g9hQzbrK+QAViq15/krQgZg1N9yod1hng1380FTaUtundLmAudemM/KkkRhR5u0Xv4rdLhVWOI
IGRH86mazGJvtsuDat/CzwrCOxiNgaj9DcUWL78Gz5z5cJ1cmSYUcTIwuEz6RlRgiblF+OskAudr
FFLZOcoxVULxCAhppTwIhj/h6xWuuqwzFWPNXE9JB/rbPBzbkzhR2Mv84ETD0V7arbcBIEGL+bga
b5Dl9AyJEnHCLnPM7KuRlrSShiVtIQg+TengvOOGGvkdbOju9jsbHbVVokZxLK95hGK+3dshLv6L
JTGRgWOiaJrvCvZCPhUaVDR6Vor4r6b1Zq29GZEFSatxs1KHGSgDo5UMQhPzn8GGqTDgPfHs8Ezo
8LwZKYcomegVO5GKuOnt15c+/ADYs7eQBHnYwHkvuZ8yRT6qQFZU+/mhaks/5JeDgJBTFBVx1yd9
WDPan0Jx47uzlR4hdH99ZZLSvDaPUcqdlLfQHTnh2DhyI4cRZMSy8WJQS9jFPEmt6ZmTVAhW6lUc
Xus+GmCpE8KS6myN+wbQEAIONvJqzGVrDii6mAPC1lFjrd5xHkgvFD7m2+WAlmH+Nw25j20+d6mg
KesfdMpbRLZpO+OOGPQ9g7bIK4lNH7T/H+A8T3zBiI9nNoKfgQ1lzxmxOx8k1rTEEJ9+KQJrgzgY
wMb1mUhlq9uW6QTTH2YcT1wuu8TVJMl+MXHmPjs+muV7IwwY7TZAnWbl2cuunEAjVV8RSXdG+/in
f5fzyBpQI/mbi9zzxy+Y6qHwkBDrmCtMLCkegBqLZJalR4lIvLt/t4hOiyzX57ysa+7aLpd2shi5
sMfgi/RHmJ3P1hFaB6mAqwS8w6G6nTuSZKPpYAJod9Zk+pzoc743sXdCNew25Fz7YZuT74jbP8za
YJkfo+vlNVDdtwBDqiOIJa13a+RfM7o/Ux8c0+F8z14bLatar74HlM8IUiltltbMgLYUhXe01TXj
ZI28vSAkj3xxE7IXAXjaU4ALrJSucoIab9rapoHIcpk1iFLnJ5Ov5Z6yiwO8Sn4tW1QFpGEa0n2h
V2zEvgaPiFKUJmdEz3qjKxdEOm7HLyMgJEBT1cNQg9ZOteGnOZto0vnI/6X8JQvvAKQ/UyKDBXr7
JVJxM3U+zLO4d45G9sapaSY3THIksYY65XtwOBZ2KiU9tUipLUjUzS0RIdiLEldClvgHqroeA7s7
FFxIozThKdQhCnpn+pXwkTzNm5XE4P4Q+HCiR1De5AwB7zjoOcWGHK82WWGCvR8bT95/C7tczIRz
Ietwr8Vpr1EaszPtP42Ohr8uofJAp4gKPjoVHZFpK0iILNP6rvZrRddRu0t0IB9KrmSNEwxIUQP1
clXoeaDzNkaSxhnRiHDrXFGv1es00iUrRQ9ndPlmErm215gZIUCBHVI1EVlHnwsjtfptFcWT3hcj
DpQNyIk1AWWJh+ylw7S62umGSfTY7zuOBJUb00Li/zp2YzWBgSDeX0u5HlyOVDHFdvaA1hSkF0yI
NP28HTmUtOV4TbNR2cun8VGzv8d2xAWBxIZC+DnLDvRA1KOXCLOXu4Alx7bSCHflKt6ETZe9+iQF
Ol9m9+QoucMiVsBN8K5I6N5g3BRjkAfBlh68PYsZVNTvxBGe1+CmLsVqRgY5C37u7CupbCi05hn1
hbo/NLPg80CfQ6T4QHv5PJxCVabowFyqDAZz111gKUnN5E3FclEBmDbJ8HkbqeFHmqulp1bG8685
xoaDpy8nb3scypifKYwwrHBozQa5ITGlpCebqPSP0nF9kvCxsJ0ZvcFHmpk/+y5NCKXB/rc/ruBf
UdCMSjcQ0V0U6sOCEuX6Al4/uQL8QPtTRdMfIaYmN0k2Al1/gZzXGcZAMT7qFYf3QErHLrlfJvXo
C/SZKht1BXClY9qxnAHOaAUQNPQaADLg9kxNs+vQsjDLuhiC6TNFvTZ4+aqRYh1aSlLEKuS8imY5
sPadmFm4Uu6M5IU4CIwnnsTZlnWD//eK57utY4yLxAGfeeqYSFNEkkszS/glDDYPZBpwx3unYIpg
2fkZR1f14OJ9PBG2fj0NajyySuua+bcnYGlWkCF2Z+sif2TVAtkyuyFIn6CTd1NQR0HBj1adP0Uz
v4Bih7N5DTTz2qhGyJ3j1MEd5OHmXgebHzt3FcSAumFT7coIg8bia18nJ2bwXBkfGx0uTogmFsBw
Hcw/MSWXpXYFodv0R/L+urdDeBojVcFeQCKHKVqTAxmZwJH9DgsviZN2viX/xGZUxxEQzOplGAr/
LwKgZsmRLNf/X4B0kOxWcTHCdUo0MZJo5arxZ2VGMoeAPRgXMkRd4dmk36pDDiKcF1QSz2iZDRAS
5B/+N5lpk+TdMLpzSr5etLH9cemu7jCyqIZ1HoiyQ5iwoMO+OsWSiyrrh1WFAT6IQUIzGrXiJGkp
KOfxHBXLkN/beLTUdKBpKpsFTmdrs4tfCGhmJv2E8CuhHMKSAKzBbWujrXAD48pmwifnbmxy/rDC
Bmy+v3A7p+nafEgKV8+fTgNrLDOTxvliCL+y+SkA8VDdqmAngemiECA5FovbjfE4dsltcVC3opxq
YmswiLvq3rDn/IpvfoZhgnRY8gsJ21qzPEA/8RrNd5YrVNvlD2xWqOzMJNyaZfOiKDq8zi97Y/kH
2RHpe+RdfAv13sQUweZuL1ZVV4e7ViPekybgQ0j5kTEoDF2g7B0qOZ9ily5DlSJtUtLnTSN9RvEu
vP5ThCMQCYud9jZkxsnCas6IxBaBXABSmcbIswA+Jq3MJA1mL6FD0dqT7W5bk5FOjBGQiyyYM2jD
L9y8VzmfRUTTCoaJZQ8npqzlQ12zOYTg4lgN9xM6l6ReVcjQHDuyJwKIHn0+qwcxNIakVJq0ZV03
Q3aU/ckc5donRMddTgyWpR9YeAJhK/7HOWws6UBAbPKN0eqpaXLuE29iHKTDvlVIYSDapqOTz5hE
ikY2XBiJHuhfVLg65m+6N9trdX0LTDJejgVFxGz/0T3FHEOygE9kFvjBGWthrSu49JVsHwueCIeF
fPGSNazkGtWoSbT+jHFdXetfyS49IDKvGgEuHnyo1BQ+8u+IQIgql4Mr3oAQ9QPAlAEZfxLCyaWv
YZffTvEI4YbEAZlGLKE9FlyugMt85oMZ9RjN0/Up6sp+7WdbIzY6zKR4hXL3I/6vaXt4Qxvy2KTq
CH8IgQh1ux3m/lbh2I6fFhiJOQcwPYOHyK6Y3uLJxY8jn9kjoH9+F8ktIKsfH6ZTdMSGLSxH7Kc9
CaJq5bDjPtHRxQFgzLdEDewxJnr4C012IKfJ+9+9ibxoCiy6Casb+/AqeK3Bkmvl47SYbIAHLAUe
nKoaPX0T/PgwD452F8zAAXmcCSflztVlQ3ZOWCemXQRvN9TRCkiUTnx7kgsUWC3zo/tpP+n3JobP
lA6hGwNfpgP8D5MbP28UkTFUCPvh3bbfm60apep4wo9LNFw0am9/F62TTlVSeKHMbpzAlfGW9fzE
WfAEwjFoVHpl5Tsrf6GfVTsqNdqwkhpAF8qZG7OaZzPUrZ3hsNiTiItWTNcwg4E6TUEwddlYZqI4
MfOLN5LoOz9zxtTkB8wsJkGI1YM6BypfoO+FC0OxUiGznpETstyuWeyl4g6X8cd2CekO6AReR1tA
eSsQ2tIjIctyZRotn8r2JVYErYCXeLRxfG8Xlv/YMsqw6PhO08f8MLj6y++8Lis+/mF/wUShHJs2
59Ihx8YvucZyZrSRaIdRv0opqq5lmS4gGW39teWEkwQU0BegJjTZ1mHZOOemClcRdG2H05GQCxL5
SOq/EOAHqPdr9QTNJhhFtU+hZf7o0gy2WM8VUqiuroAHG4FRN3KIjmhtOu4OMLfI6oR4Iv2+fE6E
8diwxJUSgy9b2NJHBiv+WZE8kxZ0yfjpT/TLTS/YU4hG5CsdbbUt1lkEvDqjayOgWreXsN/0I0Wo
4pheGJIBXNU9Ej/sWI2gL6O6VQMJeBvl2vLGW0/DlllzXcVHK4FG70n2T3VxdpIOnidPoCIfpA3m
neRLectXYX7DR5WaZcWhgV+JKigfNVv2IyZqUZytdRj8CTYhDP/nJSzKmgBpeyD2n+ajEjkPhUvO
di3Cs3Bx7BQOHPigDh3zh2/gU23nRtunk7Y2B25LrgL3RxIR2YuKF4zuqtCBMRUdKhFGbexdqkw3
e8riSWnBVM254emX5qt+u9AhID6wg322paOSVWgotqDwpjXJAiDCSXczgVrFuSwfs0dgAu7EeT5G
vS/p8OD8a7G9iBVpKuiMoxPp6ys9JvRkvbyxbk4l8IBMQp7ZsEK6jAY9CzMyyYgJFd1fxOu/F/ZY
bzWcxcqJVsBCXo69YL+7+hnAT3vIicfyC+0KM5Ybt0PjgdPQj8SZdzBDi4bhg6OI+DGDB98SLZuU
glHc7H78+4Xc5jGbjU602ab5Ov+X2aUkZ8t5YhopiSfUMb7LTh0HYSui3/geXjWOpwd4eew3yohn
P3VEQiO9g0sVJxkHJ9oWT8aPeuuRonKLimxLPgKg2gBvVmt+BVQmDthkd86FBd9VwIqT//K+0C9r
5bmdgtdaTQ51xPGGLNgcSP6+Nzn0oCZIGg2k3Qu1DlR0Fo687jCzzC+/EdZpMoV7FqgzJZtrycOh
vikFGPLpS6fkI3PKUtyK0HOkvjCZ5hVDKvO0na+f9J6QH4v7CP3WgCJW1wGxkXmYA9bVb3TpX3nr
egkMVfjmDjc3pnT3y2c6jmaADen51R7LZByfho0gzW0xk3b7sr21LYACLCM0YwwsWzEOth9iD+DK
0H9edbEzZqJtPxciDdw331tEh1lPoB8/IzFCBGYPPpjQafHxTdbMqQ0fIDI3KX8DDr860CEOO2ln
T+YL2KbLSWicM3G230ZwneCy2miZBy7c8hODgTQTdqKi/02YLZAhR+2t+eSYXHeCH4B9ZQqakwIx
eW0CHSgYTdSVlQkzuZwXR95r5iaKZH3Gerkm7O4aknbYeFp1fWL2KCzB+dVgHQhvmvh6yWwy+yKP
bDGZMywHJmBZ4xxbWW/IkjCg8qW+/FwhxsEScVo2W5+e1Ns7D7MBgaVd8L7IlknrLK3jVUEiPlBN
U1YevRLInZNOUGkkwmd827MUxIg8ZKUnksTwv4JYwh/mfUYR706g2ryNnio+WufDmRn8YvikM232
h60G4D3yK5oH97DYb6dBpR2dM64UEjTZJ2tntAA/kY70awO8moPf7baFdbpIqwWTII1aLWvcWBgB
viwVddwqsUlskrHVjbWnjBeW9HE4FVt8kNVRCJ27pzZvCn0DNEpUf20FWoojUouDp+MemkaowBdN
jWPebhs5UpaqSv4RNH+ewo/12MbYcqvX6CCOJ7m6p0XiJf52Ua/YYmxJWTnSApUXHdKEACqmHluq
KZR0RmccW06ZOnf36HJ+z8woTrL9yuVdpdgtZhyp3/Lm5rLXNk5WPtXZhejQwEeHqPVX8+L26B5t
gUTs9vQNCA9qOdbnbCXctOArkghO+MCSRkSap0h/dYTXp7yb5ksD77Q+0rzn9OVugV60d5YJeu4R
RVWeWZIKceaIh2SLGj7FvQeniXOmVbChI6C4bWiPfzYNTDfhxJd02qawENPO7wanNkt2q/hXuCRO
IQzaTZxERFj6OjXSQrNBSDPducnJpG2GS2v7qDXQOiDEFmOIkmcZ2f5SoQZR45gOxDinPvEbxklo
ezxctd+q0Nk/BjGWTxKq4vrQmU9iOGvLAIiQtsC1bWeKf3Tnv/NxtLeNR9AFRkSKFUkFUelwqC4w
E9XEf3enW3y/vEqETojEl+rPdFGL1Uv8T0pmLPlHsUqquTds7cOijkyX1lVDOtHUADJHtpbRA/mR
x4hzWtqcfwVR5qTJm2LWxuUorA0u6JWo47TobkZ4lp+rB6svoLiknmLAyiVdhDXY349FZYA4hyXC
vuopEOE62u0tIrFxOoBQ5NmeP/UaSDSm4dvE00NW63K3r2NUvo6cIYE/uqEjJ7cte1EsgwAc6qsj
dqV0eClTHKoldxqMFdtM7WYXObs9QqkWSKr/Gfg19VvoCt5lDTVw1tG/zTyYspYTCf7+160x4cHd
FWb12edgKtTSDrZ5S83b1Or/GX+/XUzhuK+jCoCmG+4CbbxWC8L2urHkbaPfSB2ZWN8MYu0mhYGE
770qOhc9+u076+7qUVEyXZdyMZjo9lKeVhPMk/XiDbLNaPBxXaYWx9ZvHj08Oih2MY11jHCcaUC7
XsNL43jJXlUhPg938Kc1BJRhgGInyvFFPXUQzk7sqA8dZdLh9GziWOq941g+sYIiBO6KSnRrAEbW
DCgguerFR3ehIOgCBZlVK9+SpE5Ahl6KrdYRaPbL4cX9F4+Vl6MTu/ePpyPTa9+ySzc1fV2Xvxjr
mBI4azMuPQgDOMmcT5O4uhdjX8YAF+agfEz8Nl7MpY9ZLhaMfSf5mfj0i9UR78d7AbWfPO7KpMFG
ZdN2XOCn3s0j+QEf6eyBHlgPuMvYKpjeNqrGWS57FaMykZhUXCFfRp+FrjBg54sSxZO/+KRSri++
gBTRS3B+rakHlJJ0cZWxA035HV1+bsFPOtWyzsg3dG8FF0cMc9093Drt6XSBHSn07HyCBoZdm/Sm
Zs3GCVDyxq+Xna94uMzxrK/HDRTzij80fyQNu7C8Lv0M1S6SY6FrXZc/HYXVM3DLC7NBmL/d8RL5
pCDqP9h+GeCHTGkExWNO9wdlIYYilVjahp/m5IlgE4XjEvGCuXDy5/+p7mDe99ykGL3TSnUBx6Zo
YCObjXrDMYL8wZzM0iBLur4xaCsvg2eST1CLUyichE8+vd+eZSLSHL6mIX9XxFWQQG3LwA8X29Hf
uUKBFyjfzOIa6uiX/pm7qDGSbqN3CxBB4MUvWDxMeIwwMdBVuWLhtM2c4JDIWP7ux0Z2fcDySAdC
YgRUsk7aQa0gHEkTEU++WzpomsVo+QUNTZoHXl1aiRGN42ohrGdMTJp3c9qIK6rY9LIoXowoEGRT
ptkxIHNWf+PcKotJELDCHMEpn1vDYHJsA4FPxXhvuX26YAoW0ILF0iu2uV2HXE1pDuKLWNVFcfuf
Lbe2mfvrpILet3WF1DCNVSeT06GbsSAZI88Ca+GVC/TFueVWp7zngsnyIv0WcGltIv9KUudNZZs2
2rI2Fknk3TpWprCUX96GOPKfCxX7B6Xk43PoVM3FG3DYTECZG+ko+4ObdQaf4rejdTIKcWg+GXnW
YQDyCF2fI0lBBK/uF9urwqwOarBHeabTApST3uEGIPzgRFtRukxAD7XGdrHniYTB8yVj5jAeIMcm
HkctBoqXWGGjFx6oTDRDKhHGcIKixHUpgbhRlTf7byuHmY8jL1hQrI16p363wUVEXSqu1ZYJIf6+
Dlhst1UR5Vpd0TVsoSrfqCJgbTt1sA+Y4mdK2zwhqs0XdZyE2Ga2L9A+SbsYJC+DluidUcVf9Xcn
KoPpdWUF9mHyUMdQfTP+GEZNMDSTBOQyBXnx3dE80X0o+wwi9NBEaGRcdlFihkISYAud9z7HZfrV
4XTsvxGi7fWdTVJXk/yXEBkHqeLDT3TSNAH58V8la2AdH1w2rSbYxrDIT9BQasY7b/F6YBIoiOxl
PVhrBZ7j8Is8fA+0e9NGXD3Ce33P7PRymFJw2ZgV6xrmBf63wvAjuu9++2/r5+2F9jKms9/mdAEa
7z5/R3gZXGXB1WOtP8JycY59840o5HPrnwspWFTcNbzATDw1qGqG+QfvfWTHcAScF1H5oKq/SMa9
ufYlh3khkBY/EoC2mhGQ5MJhBKRH/bchEDvEeCwUU4RGiJ8aQahBYE0jq9r9+IbZP4IGWF5CbPl7
1qdTpIUdCWwKpmbIszEjBueISvtimyWee29ySblNG0das6fuCmOAk9h66VbsomTrNiK66ynVDBdI
VZ0GmhZc+RME8+StavhPy88I7ZA3KSwKIut1RfKCDrrJ2CHLWrVHkhJ59jVPk/rsQMXd5oKIBzBo
nAerRIhClvCZVhwo0HtqCOY+vLlIOojxEWOojK4dYjQj6wqQlDxF84j4w4zfbJ4XhjkhsaLradsz
w46xJm4T+VNatA6oN+ABKiJgksyMQ22gvtjVe5iYA+eg58FHew9VG8AaGMjN5IsncV45bpID6/Hq
3wioVQ6buHXLuc+brSxglzDMId3IiI/zO2KxHpIL4HA4gYEfirZ4UpkPWYRiOyT+5c8MzCPjdD8e
1StrFmronhohDCGdCzaJeIKW2DzgDcmtiz1nM2ajMhFaSD14rkM=
`protect end_protected
