`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Y9HJRxBaEcwy43nSU/eJV60kPFuohObVG0NM1S7I5V/ohZNNGfbPcbco5t8L7B8ErR5IxNvKTHu1
EtXiLSKyyw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ikzXuOXdd1YkE5w51T3LEfzPDCseXNYFskQrZ9725xIz3i+QRBENpl2YVsV6ifXcvyeNn9CFrXCb
Oqm5MZgtIlL2vE+FGkaVbZtqoML16AuL3QtsWGCoalsP/VBZyq6BZCV7GbfOebCWmmRqsu8E5LFC
Vz+42aRgKBUqMzv+33w=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Wop8QCZXsyrRVjkXfocX1rSG0Pkefz7FSlt9AH1pz0oQmGD0v/seFy8/WFvNhuPXhMbN03jDz3f5
cxHGZVLLBDbqNXa0cdng7wb/mpTfHwYl2or/AXZWDp5hNQGld335iNgMDR+wnVoBnsm1PhClrZnk
gfREa2cBhqNzWJhpvkRdpfiax7U0IngaAsR1SE6/5aNFJx4AWVV0slvPtYEXxEQYNxDinMOLNqBO
7M1qUiBdx3g1J3PF6qIiusstHgSunwr3ayduyjH2PCTT78ZvcvOezd4PJXNq6ol44kwMLxDzCiKD
aPH1xuriuGa6XZ0Yf8vqckM192EfBzdRubSJfQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sVBph8jSA4U0m+NJcnjNZLz1cs3tB1pngfWSb58h4ZYHR4p+x8qv/+h+zrYs4GjtaaNwRDe7I8wC
LykbBzNnefUs5OL4AfpfuwiBZFA9NtXAp8pq4vNr0TInG0olXyG1LAQZfINapt9UWWZEyOHI/5Lz
4zkoRFOv8uMwOnx0haI=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jtCigJRKcuRDsUxXlevVyZHBhqvlWpbiZ2uObbPNoydyXKLWDGMKVXOpqYZ2xnt+jiMgPnzRdqVS
b1zNPeDZKvy6PZxfL6kGBRouiPUv0l3cbMViJUO4EdgZpp3+vx3MCpuUpJ8r6xvC5eiaBLlYHNXX
03VX4gcvvxlBjzpFE5pz8nWhzo9e7xNthfIWzDc8NARyi90TR9eDgwE8b966jNk07HzyAIiHFitA
Av3qxobNdHv4q/KgXCeb0uP7P2Y+8Btw/Tof41b/KlrVF4ic9MZzxRNkDXC4wU/X2UpKJcpfHOki
3jEMifY5UR4xnf93ujXT7ngpdIqnzl/TNwogUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4832)
`protect data_block
Q0ewdAf5wH95WFCg3LntEtRj0ngI9Kk7XUe8Pc7PTuI0WRHdTGwk2ftW5uydtOhqbBJlTSToJegH
Ed3O+h/LGLHAb6udZ6a/U3AOyFGsqq12Uv1oTqGdF9UXMLBaCuiXG/fK6XhrEcnvCe68rkovdIDf
d4aZ3pStXbDDtwOEOA+eFV/5JG7n5VR/021R17IoTMPWVnmRtVI5tjOpNynBjuWHVDjnY9d66fvd
VT65hq/o2bxVP9R/q4NqOu4KnKmWE9zH1j9qSdiuQuYfZmvfJHGOiK1oYSKz5w6pT1tWFf+T7j4b
8rJhNMUQ0ghGfgiwjBOkFzB1TWAGtGiZsnfC4jCTd3kXnZrg/B0krQzMQvVAxGY4MzszC+VOFfs7
ri4vPrCfHwbeuUw6/uZJaxf1R5Yq6GfrVmQgVItTDfCU7okkaiatG9ikWO/WXNDTz9R6nfBuRZ5O
NCr8QhewM5xZI6dt4IZufEcJFylja0925QEmZiJr5rC/aZVu0TwhvJD31t0G2626m2eMJ1zq/Tia
87S0yRIx9QNnjKcNkdO1CG1LC9Et9ZvDO5Vhu5jQAZ9pX/TkfHJAsWSF396Rl8yFVhAQI0fu0qSV
AwMZ27Nxh0h84BknrR1XqAKFn7GQLTl0TUShXy5JGoATgyccmxtoxbIsefbpUgz9FqCszZJ7SiQS
Gu0mYW4RfjjUlb4IQNiXECiT1ar3uASVnbnDsZNht/HR6Hmw9eBwpzdQ/Is955a3/iKYuPsx+eWF
AHVWWNm5Gz75dXHzpLJkv3R70GwTrPuBbDVCev08l2Hff59PvgKqmjykSTzAKiooyyqGLwALcGx1
Ygn9lnZ2y0HdM+bjoXF7lHrZFU2YQtJJXXMfmYiIRdfW4/ChPfkPEHfEklGOHA6OtXDNY7Vi+zJK
5/yCGDtfG2X5wnDIS/MY3yjPWLPJ7eIQJ6pPTTSYLPOyxfGMY2ZKKXZJuqz1lr/IB75toHCV1hEk
1KaEcETtfEz8Voq6RfSk+wzcWjU3viS6rGuQwEkpojMz/RCrLLqz+QFMRy+o0c+6xc1rkscgrxA2
mlesRbAXSP3SEOyY7rG6mm7qXM82BnfQOSMs3VrfspPxSCotSs5np0wJLYlUaNvc1CKbBKap5qCi
PGLn6/EI6o3avhIB1RMmIU/sqyaD5BKclovSddejral3QfifVKfuwgUUmkoazOoAOlku840PKOVH
jhXuFBjHHU5tyP7JmRg4JZCNKrlhQ+Yh+l8cMapcKK5MrHTPYKfKH/xPidbhqACkI/Q2vmAkxapw
+T5wCJs3IlzXhu9GGK5bnHfU6UUxj3ELWpg9vhY7/5Ge5H3aTM75ECvADcF41JGHkbvjBRhXCVQo
L4bsV4Nb3eeERSXRoGW3+PSX7q7OVHp6nLH0dJA6UPhsm7VMFVN1rWOh1WrUHkYZJTjOjQQr3N9B
Wha/7yQP+w5t7sxLJjnO0VX9Kf/KzrLskplwyhki1WIptYfbXfM+6vUOYy3DFu98Jk/hfxN7/j2N
S1J1ni73a7eiOae/zgxqkX0aXGLioSMQDNAKBALZ/PRt5WE/rzfUghvTO6pUzv8gtH3vZoMfsVx5
aRXkwziJSsVNc6GAVyTTy8AZmCOd3Sy9ujikgdG5LYRBLK2/hHjPxUI53cTRGwFYKmzNI54+mGDe
PaR46LujlLLCCGffN4XO+yNodIJvSjqgBJhQho9C/PROjvQPltBEepD32BT5J2SkvZOMnWvuhCA+
Dt82XIYwLa6FEJrRe42qXm6BKpwQTmDJfultChrO5NYPm12YLdx3G+dkUkGvm4WrpFM2/tCj2Yqx
bVgvddgemlw8/RH9pbrKJis4dwwzKuCvCZ+v7Gg3P4r5x+bVm/beOxHnoDYJRP9+1+Ha0ot863Dh
hudYpr5cxYmeI4Ya+0iTvlyxqipVyH0L0VOkLwwK6+/3p7TRF1aXKEWwGdmUe9VqJtIIZ8BQqKVD
Nz0XFtMqMvQe5pEy8H5oTn//jvTUv0B+welBIuZjfvgE/nncdUbFjRGazl7CZ54je7EsjZN4OeL4
e4EALCjBr/z6EBWJOdidSMrFmF5zWIS1xRBOEdYAjARQeaAjPfYz55pIZO6Vi+LmrwlY7RtY4To5
g9Ko3lycNcUC5JK24jnOuNDZeOD+RWWRiZPH5xCi6+URulMOMw16krpRaAw8Y3dJ06omhEKZRvex
M8VpAgvuKI3LIcg2+e/d7uXsAwUycqcN5MI4wdzKVsmuhK5nXoeAvM5tusiNGfzMILvXoQInSjm2
6Wne4mDeIdUA0n6tJntkOtlJLwaTXjh9hXlbQQ7qm0ULz93iWpl2BSHQ4CyDE8YUKm8JIbn0Ny2E
wHKBwTrXCFL75ahfwncULNcEEjNPLdDAzKsPAcEnCOqhHfP7DLpS1ENbPVeSnLyAAbdu+2Ff13Do
GxX98RXaNXlPhoWFJ+l3x7cPk9yNCCMCt49rs/YrQFFf1bUxN4UP1kIg3Z1+mE7d+L64omMzse2M
aPfnHKNRh6oRI1EUFcgIrQxn0xgixCmMePHm4wSrCec0HYvoGyy+LIV7FEFmxE7f/wzMIRC1cPIV
XzMlccPiUlIHrHey6azdne3UP2AhonDatrYT2THdG6H/hDA2JevxvYIXnRmNJ2vyxsME0uMHQZ6p
BsaRi9dkpAGg3DJJyC6XVZk5ns7nQ5tdNM2H06B+hC5svym212pC13rfc0cf1HK+HGze2Sphkkl4
BQZbu8KsbNdPuatTTOuret5evv9EKQORkHMZY2ImnQvsPI+d6MDHUFtkZGIrQV0Mt37hWeYLeToy
hiJ9OQODdHShxibliKibEgaL/nRN8aRjU4QjFIF5kgKGB0o5xQzbEw3qQOetZcv0GqQuth8v5n6e
27Xt+3E1nW98IX6T1x8K8ypmNfLC/UYtmj+SCULSCpnyXg4Hg5Qk3vSau3kE9y0ZTwo23RWi3x6t
wNTjdwplG4ccXzQixXtaBKShf+kiIG1VWppCorPBlNi6ofnaPsYUoVZax+r5vmQW3+W4cVPQk+18
jFhnCEVAT0FI8TTyQMV06G+FKy915msDzTGDBnO6VvXU/V01rE8Au4Wd2G4xeASe+4KS4tUm/D7R
w44Sp1Xv8zyc9B4inn6zpvbgRzcGJpLLSQAcPvHVcf6ty1ei/WGsJprBA/E8DuoUuPMq1uqgLFso
JBCjna81sTsJQ+cJf815zMJs9VPJYCIFO51m6/g82d80CZlSPHxi0jmyV/pHyf7UbzerEygfSeQZ
Za8DfcciYlJE/BWpX2ifEPL4gpZR45ZibWEU0TRb6cl1pN61rKnSXFb5C5/IEAatfcC5VO8aYU2P
OWRC/Gqwc+M28lvNa/c8L1cdbPTk1LfXrrE82MSoE+HqhSWNAHfXcyWMNreIKTUUp1oiWNyjr/UK
hTSMfOT8kQXFkz6acac5Cv9Q8QdC9FqRkry+F05MlFtxKoa6tAFt+zT6TUqECgXL99HoemjLo1v3
c7xdH+CWckItwhRwtPAFLxppA2m5eusZMpo0Ii7WNyfxNu0wFOgJW1WhiF5bPsXK1kYcLg6AREfu
RnEzlTK3OXn6wVe9cajeAsmTurvcdLPyQba4F/DRSPY041NB5t2sb90H4RFMxKjHX+8BiA0LW0Rq
Mw6lIXa4cjvFaBpKWSXd62XIakSMaI2VKE6rHhKFDz8gAyTkA4kzWXDsYKYT1/5BlEmgKmFS74BI
cZhw8VOH0/ffwqwmI0zBdnXGh/MRYl+VL81OCB7qTSqP+zHuPYmRBhCXr/EIsuxl7eTs/4HeRMrM
UNN3gQv0BTPsl/Hv6/ICHutyDxfiRAaq5XkVyoHvZC4x13iha2dC7XH5utjoVXeBnrkbxeGrWmLS
PRJsmCyi83Ki2XXuzxnz+Kuf20HamPudM7RuI+8SuEM2tDge/MCFwCKM7x8aF/cwZVAZkDfZhp6a
bC3yZt9+x7QVuiLr2xPSaqGn4BWlE3foTwq3ObPUlU+d1rwRQN8pS9YOiYB57s6nYcfl/rQLlbD5
3CnsAUzNBtgWq8tNprbE9U8rD6TVm86/eoRUeR4+lsYkrNzJqbH1AKdxWJv5dPJhSvolwq2EdvwC
w4nezkniBnV+ulXIU7s5KOHVGJKlFx+dUPy/xphSn9gER66hjEJ+YHs7XX6RYWX87nmVuFl8flwo
0yc3kecuLW0uxfXKgRGoIVRdA/tHm4QWhAf4udab11mGFrWjFWau4ZNloumv7seb+f1+rkrHS9Dg
S3A1Z3k/4ha5sdg2bba84ZjC8RPMczOAoHxZAAczWLhx7bWdf95NohsOnMaQBKkuKPuROB7Zr27z
zsaHE8bmJV7O118NQEntW46TYDR1Ytf8wsFgRFsR8MFBsVK479gnp4MyGexas7h3ufNSHIL3nymp
a/4WwnRCYRPGnip3QogH5P91hyddtWN0jY+eCrIR7t91o0xbKVP0xO4F1zO+auPmoLINZAKuD6K4
u8rpdEYeoiNmAp/WKPypoqSiIjz1A+toiNKjJ2JO84r5yuotZZOVt1x26ytUHjsFmjk0X2wT5m1a
4AbsFdimYLIag6ZqFvvv+peBnOrAPzXgVGgynhk/BrnOaTTwVCYm+G+xUXsXcsJVYwuj3HFpgom2
UBpTUcA6ZROCZ7fVmgz5KpeOTuMC9CxveuV1fjqk7CgYfQpFfPUE4t4lxQHsiodaeSfRYjzWkbJ8
CUeWckp9LOs6RjViqJJV4MCkqUuBrC5cGhH01qwco/Cg+aseig3Gxg++jfr+esBHtujJenkuEmts
jn6XAfYhl2U+VTVJcURy/47WHAVeAjmxht/1sYXfOycp+OmrmIDRZ6v8uZXFUciZ9mOqq4UrxKIi
J49+cKLeREeZhBs4efN/cZfsceUmPHVl0xPm9TFC6a8SNqK/RmqUCzWDOBxqhQPeoj04ZGExvJLq
exwSkex0KTQeY8fDzLhmaZ3VyOe/vZ4wF0xZa1LiQ/Mt07cO8HIZjHQs9CVgHSndEm8ZHAeJFi23
tOSqV1YVSBa+oLIBLJLIZ+Q9Be92iPR24DKAUXuf32WKXlgg+YMMeukiNWIUdOLuzZTBqSsYXEQy
WT/YsyTnrYm+OC0yOti8qflvZ12fv+rXc0Q264JuEI3mRbvPosU5+OULjTxT4csEYO2ZEtWNyyrz
GgjKqE7kqm2Kr+x44kiWHbcW84W3EzkyQE1BIj8pkiiHlbkr1mp9eYJFBv14HmcrDDzce9cZzC7l
77S5H66p9ta7KWtAVssQGvRBAx+xaJFKXvTX3vlZF4f/1RHEOEJbOvTNY2fxWbcacoTTjS0ALMvY
HhUWbGkMuvMfRKZLyteI5+BwvvqewNccq012igMyo4BgxA5xEoixZjM1ngETZROkUBn0vAtYzcNq
HutWm48Di8rP6162m7cxKGK4RE9CXZMS+C4LLqNT4f5/EIUvr1QHeP2UonTAlv7TGcqM1wwPZTjA
UAidYuVyOtEYa7OBZnRe8Yc8gMtalEuH7vy8LPTL7F6Xxu/7DTdwq2gEUBMFDG+Lg/MCGHb+6iYe
aD58pAZkB+4KQXGNc8oHc4hH9CzMNdD5hMoXXBGVpORN9QmEspyKNKIkgICDWpMyQppEgUxVYCmv
PHPozOLFVEbcL9RN/KTprki+cZIHHJHHg+NXSFLGeHMXroIxFMGlpF8FzcIG/ERe/z1lzZ4rwb7F
Ijk2683aW6q9V+R4SXNjxiiLQ2QNWKwPS7hdqHxeTfj9enu/pLPaTQSDmEfJ/iBLqHk4bU18SloP
MR/j+DRgfC6NB4I6H4Cb5fKtlyv7U2uoEg49/EJHmSvknHN6nj1YR793daNnCwHU760RQ6yWNFVM
maYgwyzeZzsxGZn7yccGxe0U0WmuygSVaHJ0EcMtdhh921YvUufghqcxwXtLz8GviJj2e621xn7N
r4iufqNiGRIMNOnbx1+PykS9s6OGqfIdG3fez/kyCSG7N7ARjD9pIv0yYNhFEPhaF/nB+ykb2l9a
BtkOM+AmiBM3PE3nT7uGa/34s+uA0wt0lhB8MudeJGbqE+cIpH394kU1yC4C+6EalnLWAL8OlBIo
5xlt7+fP60qZQpndl4/3QdZk/63xh24QgNi1PKT4cftZzHBugq/kkSr80LZUqFYDwVDNfm7d7t02
3m9FlKhoqyJmJyESsGUDPaDVJ8+Nfa09Knfnn+77Mi51mQN6tdzddy18VL9E3rXO1GoVYnJCg2+p
4oTSlGwSD4GMGhngtmzMlXM0zAw2GK1blxteBQzI4WQgKHv30gU5Yb5Q3P/s4B2/gT8ZltTPT48L
G8EHm2pHzRi2UsnkrH3O7ojqv4s/7bngE2AhLmvQqR3/eEbGh7sEGTIXhMGpqqEhyYip1PaV8baf
f6d72h5+bGTtpLf/RBzcDdBEPqRnZ1dtXJJgjPGfm0sd7eqiY5qnRcR5eqw=
`protect end_protected
