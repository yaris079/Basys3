`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
OgS4ZWdOBzSZPVDqqnHcubrvg+w6I9QnZY/XYS85W1Wlf86f+HAY1yn0j+OGYxsVN24/31l6VAhX
5pnR6YIJJw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KBCTHljGJPJnr8fV/hhnc5DoHM01gQk8zMMEnL7sc0rJLu7tIeRJ2WyeNjtdWwoh0vVIJAZqwNnj
J+u5FZgHUg+VBNE89cCUx2grqy7ksEs4E9uogRjzQZ/z4wwtbfD/xBd4+DM7SNQ6WYvRwo5AzV4F
mpIhuJJ5A7m3bU/KyLo=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U4UougvDjs8Pi4Fhu8qKkryE1WNDBT2FJZEbwkZJBXJ8CvGBtRBR30cGpceSbMmQDjJAyycYz8KD
PIdB5jPQhPz6E+WLWxD/WB1jpMFvwowi5tiMXJDpUi4ZP364T8+gd54gC/7jf4CzpOB+wgRzy1cU
ad5C0/vT7kT16tJ8gP+kurulsb3fvqTwq9INhjqZD8WbHsw06KzOIz5BnIfXJ0kmYxjgGVX9cYzj
jctKHhL+Hp6rc3RPeJ8MXdrADog8t/3EfTq2atze7niiFTtWeGghuChlNs/FF7vsXT9Lo1qP6tZQ
xx0PDGxjRWRGEzYuO0Ll+cGjlVF+h5o5X0gj9A==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
37u8HydrPsfLGwKkD5OVbbp3U/ynRZjfFikHzAR6Dvovk1XWPpjZ+gliPL2go4juUaMY6hIwFn2/
bwqFnZeiliEyIICaJSNuG33bGqHVx8MlcecQW6GiA5bxpu20K3CycanGkjufHzQGrCdBTrhxUasd
+d6uld0Y7UDDjKysYeM=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QKJ/YVe/U7mV0sRMeizuAYaZWWn4+VoWNYO3Y7FWIK7/QggDGvT6XM+SOA+OBD/+zirg/qzK+ZjD
Ym0zpxAIEpZ+UgJtmafInc5hSrGEbh0T9KjP6TRR6tNfEJBReJ0nNxHhG84xIcrVvLzlxKAhewfq
tW9dPX91Id+s/PAelfNw834WKEkn3rwymPUCaIiCpwQwGtev9hofxahoKZJm02KUu0pmCXLZIoDt
Lu+RdEWaYVFsXW34bN0H5DdymjKjZii1FcUTxNr/DptYOewi5oqHKG9DHXqDxJJU+m+M30hkDQDn
U7mZJsj60AN+VHXX7pEq5R+crWoqGevi9myQMA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13136)
`protect data_block
JYjpOh3sWNb9h/rluaobbm+Y6wLnskMO9wROarWv6M2963tnKtcby6SFit94eHxA5L/QyN/XIqES
83TXBO44CrfArcAgVdEHR4oEZnfPcE+n4sb8WSEZobYVX7fnDPG1OoOJy42X4rkbjjLiiuyjMw1V
H4BARZNI0yOf+817J80ynMqIwRttaEn0Fhhz0gEK9GN5bti6Ar+Tkee8aytlq5qGUeXWtTsMYYZs
vJJPvG/jRMT6tqFGR5Hl9wnXFDhYJ5okIeuzJ9h9jddLtFO3IbX/oSCW13QaHN/6smuKGjdh9uRQ
ynmgAwBWOp1qkoedK13eks86MVtxd8CqxyiUml9ZOTshgljD7ES2PL8Q+spU7VAkAyZmCo8Ki3dJ
ofarXny6+tzoyK1eOmPqO3vXRd/Jo0CI26YDY6VTeNei5axQkF0rTHZ4Ob2hMdD5Z57c9gnQAEyG
21HlWPNSupSn+OSHh3xD2G3/4QhUohcpIWz+cSLBm330a4ytiWzlNT0I/uINNTCouFkTvZa5KIa1
AQLVjHnzcgo4barr7zUKAk5eZb8I8ERDE/l1/tFeOOVmdg7k8UBZkyFJnRQyekdzfkr2Dc6C4JSD
ZlAuNfp0FUaanuMK5gzqtX/Hz3JjMrrXSn2l8R4VL8sbM+15v+ey1gQVmIvwTgL9So4jknuqFaJo
xZ/Ig4ZhLCRM+xyzg66+5edvJZ/ytNNrp6C1kqSfbTWb1hiNswmOxOrOvr2UoPLQXues+zYjYEmO
2PevNA3OD2jCOGoRkDuE4b9boEc+LXQ0ehrdQA9375i/knl996oRgdCC7DHyu/SXluK8TrDqe/mS
WdN4Hfl0qs+JPpvqKQP0qQ9GpopPfMwt0Qd55ZFs+xYY3ni1QNi+WmFU1fmJ0RoSQhJmD6lIqSH1
OpJH4MznYbN0oiKa7ejb/W/HST8wNpcju/8OrAFPfQ8QHYqKHF2Y250eUC0AIdOuicy2rX7wUyF4
rIFY+Epl+9bGc1pJMPx0ulbnvK6/zBx+USUk24LQ6pPyNXJA3w+xoAg/Ek3pbROcsKKfh1/9jgG0
Tex2Qa7w3oNb/04iGH5oJLkJVuGT+FfakS9PEFg3okAf3j1tNtHhTDAE3fAcku7546g2ghO9nCkj
LXQRAMuDzJGVStviepEm81sG0JtByC2zQYTQ1SO8qWKv6G2cNHbvP9OwF6LJ29sy8Q4X6/vWXVUP
ewmfmr2nuI8WV23YXrCR8COprz3DYESqmlA+JYyQnKuayuEp1B2BAUxk3+tpIO/CY19S4fjhFsLF
8mi8hgFeCNaWzOzg8msOSK4kE3gB7uxArgR3xeODqJAF5A9yA6CZVV0dVPYMsf2dafoqFBYdKs/Z
Ts1uox74l85fZKCa9x0pyUe6AeGmA10tad4CNB9KUE854Umb8dVlh+ju0xWlzfQRomFBsnb7vZHC
Fc1XWSJJYTMzHArgS/RIGzJUEzssa6CInBqSynsoNvYluSNoP0NYyFwi9giT5rE/3MKQf+1eCRei
fG9JmQwe4ahV9yNSJqybbiXreOBfjxCp6bEMwAXyZaIVsy+5nXTMd4hpAQwZZgmU7s9eDA/mvCg7
mY7wWzUjYmwrhZT+A+caXWq7tVDMmMrja0xhSzAI8DXV4PHQTT+7auV6PAk2q6M2xisbk0S7U1v4
3PZk4EewZakojmyPGniDDhqjVu8sFzDnUF79OH7Q6oHsLd6AqypYGDl+apG2FuG0yqM0CqGyVi7U
oLN/2HJQ/xbWnY8qoPHEDsAF3d40CTFJfQDvVkPc9IMRuSukAVmhY4CT0L0n6nrHJl7xfC8SLlVD
Yln14GMHPF8OXcjzog+y45gzP2IVKGi9WaC/XxpRQKfoGxLmj0B9lNVJtmsj68jMAi3vShQV6HAc
tPHBQrMA7mSDL80TnEXXKw095OgUGBpC77qWDnhXSiYcSynu1JL4T+/8NYNeAKu/5c0GJg/E6uQJ
sM1tlNejaO65g/a59WP+1bG6vL46kxtw3a2KQ25MQKEJgxnznlG3q1DxJZcOlkbHeEeiQBueuzX5
BVRteDN3sLkJfxTntE+BbMMrDYpmlK/IadBhPnuQiuj2llrQukz1wEXHBafl+DX3MtjBbfdBHOnh
33bGH9QjITAtmnJrCCgP7iVo+o56dmMw2C62TJkUL3NcyX5YWhlwR3NXr1RiJcl4T6x0HQfDpYUG
QUzIzJCWlS6ZaLiIdEj3+qnHcF5z+5yTv8JlB8ZvcB28ADktkyGsEKttAfB60Lphe2aGQlfseicS
2xBJ1Sf7UMwPI6tGjKxNzFImM0ZixgLQv7hmDH2ivRKw2Xn02WhjeAghNhldty7bJy0IcOP4+obd
eboVSaN7lp2RMwOcTsRA4m3VvkrWyX3wee07D/72G7oipCMJdlWI3b6x886mlAAL+0s8Bsxb0wq2
f3zZILv3yBkqDipHvDNUgeGusPLlThRbCEW8QxTEnBNsm4Vk+mIcS16VAcwxmxK08JLd87Ei4SdJ
wKnJWe9F7YuSy13yJ601yLN86qm+KUjLUGDMJl7E8TUerAEkxlbHoAr+WNU71a7i2SDGLc9X2say
hTgRnIEgGB6txaoIz5FLFzWnTHBGL7v1ZaersJZDp1ERjgx/ov0/4Ly+lHT1yFlx/KfmGUrHoHLT
TkZj7oXFaY0otJjWcZraCTi8Ps/Syltd5Cw9Y76MUd2k/zA8xnw5TD8MhfkXRQp0dq8fSEaT9FXR
vcE9OOjeN4PvN2H2dgeiXdwhX/LicgklLDoZOLOqLCvC0qgRAYMYMGqFF7hdUmx00gKrcIl4UAjV
Pma/KkXZWSk6v5+LapGHEkT36EUzLUAgO3sESdioYvJdou58FvHNrxit0VyzBNgzZBun+alahpSG
iPCXrfp1zeF/3vcCIpzpuhRzoXh58EvcffSmEfQCMgAm5fMS06CYtvsHkTWIyw3tyTPyPscfNcRs
8r3PgtkRPU6Ex7qYvvv9vRcWmTOkpg7FybHutDphhSOwqM2CzWVhiebqiGVZeXnMOhsD/MmO8s+/
BUHBa9oajLjEOd/tw8hnfXN7w9P71ikb36DpGgmjvdQ0W8BEI2YEIwrP5QcKTT5m1/kTQiOIpwIS
rgWaayrT35De3wUIb8XMJgYrKdecOt1qbRC+wUmA6t1ksUJWy6bM5zGy6DCYyPYrXLSAV91D2xZj
I2j1UqWSSAtwFPV6iIanV7qvYwsOjuehf6f+2VSHIdJNZ1i69yXNADjYoH6WlKXQ4a+orHLZlFe8
BNgD3p3A8Eq1hmcz1BExq7cVgPBDDgI33a3bTDf7lPg7p4s8qnuVixB3p9kumz2S6U1EX4IhdvSX
2dsLfeHpBjR1S4GAWFrTP+7TKjQ+T9eoj1Xpg5sK/XpOtIVWZr8wiauQltspJ8H6rPCyvkX/jxHg
/vEiInAh90bt2wI+I4R3bB6AgOfKeTvVnUH56obJ5Zj5iiOrpcmoMDpUcdnh+L1SEWQE1/qfhQAa
FP6Jyeaxm0WtRNazzQhJRoyVQErmHRxlHy5GO5xD4zEdTcq+Px8m0kjPtsLakuaw3rie7lvF+TQt
svDX5w1EBqhp42i84Dm0u84NvneDjoYdOErNm4oeRaD5/VanFy7nkq9HzdTEqOZn8ljaBTPLyzzy
0QyWPBmSZZ3rT272ni3IWIWow+SfsC09v6S4ea93PoVde+9Lr2A6ysJ0qYMlRh1OwGCVs8D0V2jW
9OlcqQbPiZqqVvNa82SDR4LIORovMLYBll+9YssRRhVfj/Wq9xwgdU+7d+48Ut3RR3u+BJjGc9GY
5GfHDChB9MV68yO72bPibKqyxtVUqT2mkH9bFMSSre07f2zfabyDK+1h3sP+KeOUAQdKiPFTx6k8
d33TEmQ0V8lEI/PBKktxqhKTtN8MFVXbbZuW6PwCOBYu59ngtKIEI8PE9/df1zArcoGBSMkxSIMn
beSYDUMSMN89+bUMuAC1wU9eaTc+VsLAenXawO/zf92NAbXA7TcqqZhkD8Zx1/bJXMFLJtTw+BfZ
jc2Kw5OKkfR0oNWZFDZ0Y+jGWOfKeMe8ZrmmYypGjTiE1+stJPshn9hDRaxDXocsgxclyqGlfCdU
uFnXhzXc/oZnpeDq3k7twbF3bIcvLkNKz0OVfGpUh9D0b1J3AiU4HinVzDovoNIgC5P2MJuzB8RZ
CD/ACiMiKVi21Q+MSG4rLa7N74VwvETGx9F72OUGpglbb5jx0YT1x9zRpuI/gGIX7u83H47a8T84
SZgdmGNL2OmMnlN+ZaqydjJj1uj5zwxznmQgfrcvHFmYCsWKP3y/I8S3SOYlH26REolqktrH2Wcr
yVVjmC4R0XToCHAMVBHck9VVf4qQHAS5tVo6wOP1soOwMZ8op0uGAme950YFopE0Fxad3KDxAiap
RGM3yAmwLt6N9d7+a9QaRCHs+2lev4pTJ4ofN87mSfFnRkWtt5Ku5ipwHNCPSbRro8rEHHwcnHDI
jvWdIsmkh071Imo4vbnwIo8M1yznWN2szvwNj3ySadJfFTBtG/ieaVHMkvRe4+F+jPTo5wD3Erzs
3sXQjIm/4zvrbPob8n6A1vuu6oxTtD8Y5+LqSWJUvMNNj8oBIViIl3ti0wO4aRxAJndb3evS/neF
kumGG9ha4FbQhp3iRnBe1QjIKSAn63gtZGR/ouHchMjdfhg5izeEOp6THOnOdKskHfqU6nTjnjjI
f3/s6XmVxvZeQBCLdJtDYsr1oUmlqnzu5yLqW5NNQpq+kziKACq4NXNAf24fVOAgzDylkMVmi7gu
u+blK8ZFjfGQPKjumnJanRuA+WfTniU4sUIDzMt644/ODVhJ9bF5WIA/n6RNKZuNRO+xe+hbeEMl
RIpHleBSHx3Vu10j/5zRAHpnOZY+DbhCFTuf6v+xCqOkPXYLPov9M3AO+xOTSnluh1dF5mvSxjZ4
eFW7Vcmjh25ooZrQb4VGexB471nd3/5dWyi4c2TcXyLiO2mY3boM9+r1ttDKYwOUVHCpfZ8OijIu
WpdP4ACHB2zBeTs06y57Ed+ysSFDQUp7NIPObj4/9vxY6zEfJFD0Yb00ogJKzWVJFdmO8wApeGAE
5DFL7kKgGKBJuY30eRysvejG6jFvjbAzp1D/AtrKgPKYTpvLp8dy3faehMjyCdK9GugTryGM7viO
k95u63hwa3rBArRYzZy4Dq3pgY7GgzzARy8FqbcR/7XUlRz54t3wgXJBRT+5CEExZ8yCCQXlHUF2
/BmTRgOV/f5TjFfS6vDSUxJx+xZevkEjNcbrWol4FkcWyvhiPRJOWJfyCbyaswpGPlCAdhj3gNOC
Zkxs9XLRzLtJFT8xerFp4/vs78eEeXNzkuMNzYnJqa7sAhLHBFa6UyHdscqaN0oRW+JZcXcHRSnl
GYzcFiERsQbmQMaCbK+8KsRYMLWJxalNe6LP1eWZzfyoCy4PHNbVvCn9K5OE/jsLAkDI+Lr05uiG
K3VqFY60UtC/zq/hNb1wWT2lCRFuaaia+Xuv4TQ2aQjFweXJzhfC2CNOCA6OBQc5N2+1pkcamwVW
85Hrb8agMowvyA358NPvST1FZa6y2cluny1NfP6x0zkq5qOiHknpefrTPqQT7ru8tUN8Iand05G8
8gVQ24TnYgihdHLlYT/OvIRKhkKiMxTSfQGdHRg7LYbXEr9cNwkmzjh2NXMjoHwGclp54oORK6qY
MGrPpmTHfnXfihNHmWkwrGaJsw52J7TWyAdLiZg/VxuvP1FpU80EH1j3pPErqDylpPsGzJNtOMcS
WmV5uKPfom2YIZctr+d/wTC++tNew2ZcSEHqGdxAWMFX0G/r934WPIdzybnWp3/ooDI5BMk4vS5p
+18T/R9x+t36wN4Wm+yyPt2OB/vE5LjfrmELS65RxGUT4cSBFM7E0cPsMu4ygsu0P3pFF3vEPLsz
e7AM91GJAKfAz9xY+8qWMOyJFfUaH+MMoqO/pqDyYmob3q4LZyPW5sDKcpHh3zGkXBdrRWKWTgoJ
ekZXbZ1ELi2UFxDFDhsOptGP6eDUNdCE3MZL4sBMJVgz0GcpfXEvBFcvDXTgfp/tHajKVq1LrYtK
veMnhnJfWOkFUejI85Dyc3USfylKLK/WGNskARP7aRyINBjAKuPKqKBQGAwAtOB+gP0mGkjNt4Bl
uJ7H/+fpm4JQJB7WKOEpl1ZqzFpuEbixzfzDfLGCDSEKjzBTdKY0EJroUFqFbkkFsOsI0hYhTZRP
++Qx5AEx1L8uz8gepRJgcKX+7oKX9Li0XvmVYi/r2+doBVxgvDiCo8ZXjjP32smTZsJvP2A07G8b
JbR3wIJfDsVCpRmKGrFhZ8syZ1XKiksMiy9JcaXHAgvaRxV3OfJt1/OA94fMdNtc18NP+QbV+apm
aIR+XYM2E3e6f/cG2K9PZbSsJ8NS3Hg8D05Hid50r/xiX/5NZexGoUW2dA2W+/PPo+jgBL9AMpkT
cHQBkgb9REDtgcDvNtUau13zuKCBCxhHKoSyJ8oWDDzmi2JPHPJaFuyADa7UCxqwEszahOh7xdLg
imabRDMx2VA6x40pLJns9AK4c9oEBYDL3OS1o5DxzTrgUS4BDOJG1ZN0FgQzilEMNiwrBXgG18Po
4k7ee4/shbT7unFcAoY0g5y1TiPK+X1dNEx/DwvLyLw6PAq/P8qbpzICck4SoX2zN/S3gbjJo59P
XRNrBKkRABrhZ3AgsbL8K+gxIdZC8pS5p/KcEcpMuO2A7AW7OzblPNekxuVGRj2MdUgIQ1Ep2V1G
WC4MqaX9xKnywJ8d2l3OqNalhBpyaAKsX1qfiNYa0YLiB4D/U7KfeOmzFgPxI6zrz4cDPobVRSlF
5b+ACFy3UDhWdVMKfi8E2fKghKtwi9Bt4BciUodEN+Wyp1XWW1ec8raFPeRDxIVh002or7AelGJu
gARC9w9mlXOk6KTAOSBxhJuy+epyvLyvzvQ/T0b9GCxTkptbFwBMby8veeV4ekZ6shc5eNuMU9FO
/Mk8mj07IlnOOEn7M42wrzhl/hFqNtfyTaDL8YHPaGPw3TgN7e14syYUr05cyOh46V6z+VjLzkXe
14DlCV+XDBy2YPaaeJaZzBnPIKVkHUiEa1NqOFgBjg6M9eYbfbcjB0uOomwTeX3qiGaIkDFt/05W
Tjn7JRF0cMC8WVaQRq8VtoaQ661qiXe3GdxH/xpTTSK0lr+R2u09QCV6UPB0gLqg2g2zHWcTKhye
AN7wzAXKq4dyhISHRp0jA5uWXCMPRQoykxghYDpfmINnZ9ouJJYPb5b88AikD0US+N8zQ2ylWF1l
DsrTtD1XaZ3m7mRt3qUOqsGBGxHkgAQSGQ0Tj4JIpEiVeZTEh3EaKQPDROv06HbLl/8JWvkgsJ4Q
vkvp+lKhIRvRkAMeGpFapUjYQASR2ticm7a7yU+aIk90+LNUpR1f/xTsad14lo1UzWzuTZw+uHNO
NpdB3Pk/bpCNzxqey/Cs4ncvWVNamsGYdObirB3aqX6P9r1WqFTo5ntvU+lBQ9aVHw5KVGi18Nft
CtCn8C3H4U3tJBBG5E6fnyWUTJq7diNfFD3WZpX8Y7H+/MbYnbZSjw0mXjszi+jJoToYG2qj12DF
pihfRNS93IWjeJ3l5I4EOVMtYTErnc/EAhTeLqNQMvHmCP66iTOJh2nd2Wg2ectyZS0oZfD8dEI9
3xzWZPBSjypd4w+k8YY+Phhu8FP5GZ0GiX+Q/VkQUDL0XtZqRU+PztgXtCgaMYIGOdvuwB4j1cY2
e7lFaYAKT3IBFH3G8ZWGtZVBgn/bMIgcULfELR3RfFH0N/JicXRHPUU4j7Y3m3wb1feryS5aXi6Z
UnYZbhJm0+NKv/L2zku8TcSdW2URLI4iUeIco3y7eIxxfj6F+/EotYBLhNmlrf1AihJIAaUqJljR
5rvF3MFvdOdRdRnrcxyL3N2XI5WfvY9M7W3Cou3LqQuGFa66RfYOTMQEB15loA6jEwW2eSeuwFIo
tSU8TkVyYAvIXqGR7ArlA9KDLWEc/nYiBiphe+Kzz0Mo8PtvWzGYD/Wwj3G1rjIILXQTMBVNX/ff
G9sFsVX0sCgh04P6mZv0owF0/1/TcrlZYxTPDtkg0DBnXfGoeyl2hFi0Hs6C1iQqtegKkFds9RVX
JKOzyuC/0wY1Uey84f2/4z+h0ZKeB7F7/ULamhOSmzkSp41RybXqhjdrP7IiSAnkRmkbM9/MRkwI
Ui4gkkdPxiC8ztr2q4Xk6paKK3GY3k3P/bBia3z1Yj7prnK9SpSjiw0OSC/uz3zUXx8m6/zqQ153
Z68E3APSwZogh58K3Bm4Sq9cJc4/Uzq07V6UBxW/XVaVDbeISaYAahjPcFS7yObWmnqMIuwP1jRG
rQyujPHiRQ/S9K4eI9tk3ih6+hniIam70fbCFOvtJkQiwJxJ/9yz+IRy9XKWt3U7280y5yRRSoUG
vMJ9lEoqHXHUTM5SzbBi8AvSWTa/dngQAww8bsKLYXuCzXc5CyXkbNu4EV0emdJN5UhJOng9Acmo
mTN85RmgGafb/QxEuXwz0O+2bHpq7wn/LecsNFTvt5yg4iNhM6tMiKoHcpMo+zD8p+9DT8asml/n
Tr0RX+43p4sFU2KViawXrZsfULKTUQWuUvHfKzeZsTmu4XmuO8g3P8LqQl3mF6MKt48jD+N6hY4O
6QqaupznHVjUBpqquS/264LnlVfRQGko2y/7zsn52MLK36ObRAk4wFnkufNcje/roJHyY72VMTYz
StJqn2L+IMPtGWaCy9NqH2tLw6yOY3ItD0WNXTJhGXZkwr/Op5fa2HpffH/fvlOIUY56F9Ise4WL
u2pRIoSi6sUcVaF7bDTxRBmBcIbRDx0kPIzwzdm5dhdH2/os+2NgZwrRshVS1mcsmUwxU8ppjEzB
ZGbwhOMGlwqB10AANPI2UDwp2KVyCEOsAGxvxXP5xsMcbUyCG26gHrzUQt4J/g16hKtnKio3+XFX
oWsQwGlil/xS7ytVX5ttqzRTQHi5CJ4rrip+9oLsX4OfBqFDWZSJQmgu8L13M0PZkOUL7SqcNu5l
JQ2UNj/jb6+vcpw+MWd1fOQQcc0wYzQXkAGcmxYezDuo8z3fnGRAz7v4aFZByl1fxIOQuVceEKvE
rO2OJPOpLs/CyckDSKjDJX9m44ndh7/ur9d9d6dbrkMSST9EpPB9ZsWkQ6wu35fIm+4/rhFUS1G6
gj88ups21Xq0v0TvxXTE31/49CvM+ftdhqT4AguwK5hLd+Yg67sdcSQNADGMivsFVK7F6m4ZQWcC
3mGi9NPi1L4g4lZuPzs6bxLzU1uQYbM+0I2kWMkc8WmuplxDgQYynC8lwBQN2RfZhNL0jFzPuN8b
zT50cY5HqK7SLaRdff42gpTsqAGv0MjkRfj93CIm9lcNPWVt1FJJibQ+jB8MOKlE30bk+9QhS0zX
41uWL9p6yLruewiekVh+B+UuXub2ZD21pRIc5WEc5IF1Fxv47OAiIjl/HVvDkuEOy68NMMx0n+U2
JjkpxfPoEUSJ8O2U41mV4NhNqEYmSKQfayxZlRpkIqbsMQ98Hoi5soeko0sSl0/Hpbuo6Iad7Wop
D0hg+a5cghASyW+GMOQHrSsQi4ZJK+vtJbb1BEc+yE7DvoHzixJcfeMVWvMi0KpIbxEEWTaSjAjP
r0z0lDsoTwMzY725ISur2MsCB6c2pt+J83LZZAbLdE71QFZoJqNL0nYwwwpaVpEd/4+1scOjI1A7
4Xg2aBNhKjKkxxERUWrSwjQz7rl3Wq3nJibTHHnIeDuyQIVa3XrBrOMcfinIpoY33YziIsi4x95o
F/yHtwtZHdtIIaaKL7wmmDNcOU30hxIFykR6gUzhHMK81IluRZZKJQqjQ3sjxRB9Cw9NKGwkQZhh
+c4LeHbLpQyOsEecNFTyBJSqzLAryJLYOXKMfgqwm5wrdlfFlwqmiH7n7g0JpS/qq96nbIrl23tq
wYrtmXagNyncTNC4ilH0dkQH2N4rIWQOjA+4DmDdbRr57YQe1RSBynSfjph2VwEDqKOlXiVElIEt
3IGoDkCWkrULTkKzFQ27mSRYuIL1nsCPVvGnKIaJXVOyEua1/w5+oLdpi4MyCg/Bjx2DqNQr0lo6
C7UaMw/bsojkb+q2s3EyPvH91tvITGNqXg7DSw6f/5FOkdtj93NrOdD48IKsLjFj+6/4igw4FBZe
SpuPGzOUyQRPcIMxIm6xfSzZ4JteOB3X6YsVasMNjP8pONcwu7ULcbK7AY8WnEE/2jLkunRxrAuo
1hxq034spc/+LujBAHGUftJMCT002gbyms7aovClyHEu1YDiWBEDfMHALJM2PA9n496XY8mj7WVc
Y3kiPDzLu9UiHWDoaItOsd1p0hRT5MoLrC23l+lI64KFrC3yGR4VXdm7MUaCzFjO4qUzBj6HLRN0
mYds2TubjI1cTW7PviIIHQidx4WSHYetiRBddDTwZTjdg5iHFhZnH5TUXmLGuxBrYXz1/zYruYpr
GLayfIwtHsknRgdyogs3DfOMf6T4N3tRtEomvJbeiNq9cS4lPeetoBjnuoIF9iTn0LqJOhe3DVdm
QHSkx6oBegn3yR4bWjB4ygo/n18/Qf93GAqK35pw40qRfKlDay9GND1V4RlqHcHtG0B+bjmxQMRg
eGJtxZCg8sx/V6oyTqLw9w5Jxu5Y+8n6FeCzDGU/1U2hbUkCWVtzhwuWlFKbl6HrHwHFISG+Ry6K
P2Gth2VZjTvdAsaQQ9v8Co4NYOUtwuBsBWdVyfwT5yfqGRwfp/7IOjUQYhzLoiIijVH64201waAg
0v5vzcWgQNbhhV/5wB+l2NrkMh5D6r5i8jNqa59lhGpqwZwEUOuaJ7SVUi6+9MPx/G1vW8ZAOcGX
Dj4UdIWqG6Nl7cMd85UvX+80hW/s+YRb7RPAfn4ymNZsth/mbIQoUe+aVpuomhjF7GL8bf2x2xEO
fM6MCVgLthN9dYxiGqw7kvJZ2BsBG8u25x7WKzGv7fKKhFM8pK4n/F/AMWn64Hro4hEyRfi2hrFl
R1IibQb0ha7sv3YRFVgPVeMUCR6y6TO7QBOa5eQ/DvkSxBOiKOcdVRG7jnsNFaV11+KI+9lcUu+k
p2vJ1nUTWiuazv4v2LqLSb0HsP/Nsx015MeZvvsBbWA4xSsPLR5IpiuXqlTAIvR0e73fZnbTDZ3F
G7YaYtCyh41hS7MCVMx5wl0wfZIIgqhZ0yzkTLkKNAh4NQPgUf69LL8xOWpUaVCZdYMJxIT47nkP
Ty3FHECy85DcxWPhz5/oOIQaEgpDz0NTL80sfQaiMjFUFectLYHQepaC0KCW4N1tPsitSM3PW9PV
PNJVfLqvij3QGQWc3b47F9XtIUlmulwkkw6cnA3c1Nk5vZsEYG2oDUrZpk1VMD/Le3DbcYwUJ5Cw
CWya6DY+88liQk6AglxYBl+n3pvUWlXUP7Q2alYRNe1WzUFE3Q5x/odhEMzedDK57u0Y/44djILB
AcXVBgr4xKU30sMBdmDylr9v8IspBnME82zkwatkbPh4Vi9FAZkDi2i3w4T53DzA9YhtJItPt5Xz
Bmc67Bc0Bkod7fCF0T1Q8VFgNMCNkbwQDaQGbJmQFAXdo8Gc5iNadkTnWAnHPswbHhQHJSRj+aR2
VdC0tEazXt+IFlFPb+u5xaAKZuKa4ywsIUtJ/a5x7ASPJC+WgR5JFJsApWEj944x7EXbwDBhUeLu
cEwm+aPSNAaO8UIrS+700eWTt4lDkFUknDznPUuT3COZOUeqkNwgTcCFyv7O4nqdL0/d60OxW1lb
zyR9WIMzft78eCcP5QMFxscVlpJk7o1XEj5c1wnDqpwrGT6ciTZ5+p+CuePI0PTGlMngQx2Ze0Rp
h3qFlYEwDiXjyYu/uTjZq5B++wo+ShyFTm5d3oIdtRdIaB7ochOsMkAWA7Gh40i9Ldv56oDwTfnj
lilUHJrsJDmzIEY1qjybOeYiWmw1rU9kDposGzZxXM1ZP++fNSALthDRWMbAiEJFfbyTKqNYpj6C
xM9R3AVVeZrrUfDBoGD2hgJa6kCzvomNGtOmd4poA5W3A9NsyxEOlVmHXi+U822q6d6lMfHDsNOb
NYoU9HhVLNUcewkCDcZi9c1ZxRlYPGreEGjAOnycjahGH+r4B8pXU+SpPho8YbMibPnuM2h9JU0y
XgCk4mkGYZBxkLSkA3mCcNncyh4VE0Eo98l9U/XKxbHDhRJv+mlQwEkwYzqB7VYLnfhPnb+6GF6a
4Z6b5HYcBcUTVFHXrVBOgpxXIY4DCEKiJTepLc09TOnNNlxxytEBxwfQu1tITdwofZfhBmmYcCHO
XtxKqG8U2vqAQXqTUDSCrHNbupv+8QuFctCLIXNnfNkuSLqPXHsygkSo5EN6k+c7Vt+0CGDCE/yG
iGIATZPJ0VCRaKQVDnqE09QJ9/8WZBS2wPmHBeITLaovVCrUgUW8peI1h3HhuhRE6Hrx1ElEWvVW
79AqaceSOs/+IPLkiGnR4SyTdTjGG1G+fkFzmKPmSy/CwkU78u+FLtk/8mpORt+k78qITRpaJZuw
YLXamrN+x4qW1qOooGXVrkVlj7KbiX4UsgUaop8QKlPpWpiydlF0RlG5qo2cH1tLkgBuCUPSZQwU
1MaUj3iUNP8vkCcPzRezBnjD1DhKXDg4q0ilPYmct0mHMbBilUTFEZ/ECb4F9yJJx2rsL5tG1Ue5
4z5pKwg4GuI2BHQNgmYAa+H5qhs5kQA371qxTpIunWegMlk6VGIu9C1GYygarQpHHclvQ2TC7tkA
KXPR72xcI+kP5IYWeHQngAboHwKeGjhSek1pJZA8X69k9rhWwbVZmCiIwt+2SX6JuRHGZBs00txL
Uqjdvs0VzTTMOrBR+yDJXFPU5xiJ/gDxfcPGONtQ8b0PxEkeL6W2hJcq4hPkwmYbCzNIk7Unsrcw
p1U1iFN3n2iDe7NZc1/JL8OocQesrUGHLYdhTbID7KsR9QUKK/bA2TWXOMU2X6zQmDFo2M0dwfub
r7N7Vw4BaPRRejryXNZcRoaS+6FIsCNN37yEgLWu2dm8z5akprAR1tiGlOBf63E2wZX5AGZ+E3WF
t4fwJ8PjaEy3ROlk9CvjvVZelPfsGG/H/0ihjifZ7XZUky8oLbOqGbkDRN7AKQacWWQQUSEjzGn2
XxuxGL1k+jJ7oL5V6/tipTPvUaBYpXoAEXZFA70Ktk+rZRjeONIKgRnaT9Ttif4av0gFOGwH+Sdn
Fq5O+kUBpQ8XCOH/lDNb/8be59qGbEwyQqFurbVR54aS4MLfzEYrNj61GvLjUesYo3muKncYCb/v
3GC7b4obXqcMgx3qwimhCgZToG0bNp1I6oW8sRJ7/wA/8SKXLsL/8e4RUnqBrFhTJ0yYcUxvb88C
pnkLata5rjGvUNY/DkvEOJ3qnAd2pOmlxuzyodoJgAZQ3STMpzFA82/8qNbPnuUMfvO1Dp6vsYDr
UBLG8/LgiVQYovoPIBQYHunPfkm+/yxRQ+4MtQa0bu5lTzPZrCuNUIe2sEDKCy5W10YlsGFx5rst
qXAML41vZBBC9BwGBJO4nLLLtmj7aPRb8TLhU7g7xTdS7AciQ3ho1A+Ob9bzMUxABXYCxMvw1zYp
mYZ6jDyR53H2Vl4rjPsAU000bzoCSIUgkbNa8dn3PoeOM4qez9qFRYg6tKEVUUbEqGzdAvwaABJ8
sz7oEpLz10qIGQluuRn7cOhy9Vyxr34p+AA7FAp7dZwBHfNcFVv2RL2GqjVvwz0LmalprcfJb4MR
vsA8G/9F6y7izELH60baZvxgPd2qWqnxFF5gQi8h0qX4AwMureRjz2fh8AkoXR/e3oX2/aQDEhY6
KLTxjm5oqXrNE/8xtOvxrEyVEl2XZ9Xq0BzmWYBxeI7DDv8AqyCcuaHDfcYF3V6w2llRyN10/mnF
+dxq7SN6rbCy89Aa0Cul94wgycR60T+gDKsv5EZRhx443Dm/ZhmJd6ct3lHD8r+eOj+4a5LDgnSQ
aL9Ldo7Ka4x9FXRQEl7+2WdW+OQlc7pKr1R0GKFT502a2wjRkrKZSIuz1kCN4G1ns7c6Q4z6BjNu
zsav1RU/asHH/nbZedMGxlZYvHzRarkOhHG16aqY/UD+5ZMuT8bDOi8WOvaJtWnfiK+ZbvT1wr1O
vINbe/smeiZK8M9C0Ged9FOmWW2OQ+sA1N/Dl0pB8vtLrXedReLUN2N6hh/0mB0Os1YzvgmKM3gK
fejC15pY/cZkx6jLutZ+ImrW/XLcR1/3kU0FyGiX9f4UaMuPXHj9begfBgbtPPL1Y9lEyr4iiGZ7
llW+Cw1KiAzsRigeRyhpAtpZXLt8FhVupqprmliuynVZ7mpycckD9fR2QtP/RQWBtxa0wDF+HXqE
CXFLP+SqqlzZ3ytAEAGz5lAeKPpf4/2yAuG+Zh+VRFpLbQf3+fmtbggoHYbBw8Qgaw8fFepB0IhP
G1ilSqWf/De25UxrAoJ3oQQ+ER76pHAyxeVdrWVgxcDauVFzxSuKlaj9A2gzWFAs6ubCel06Lanb
1apphLYMmN4FArCJ3piBRv6jPerEBd4WR0/hkOVPbruS6FmrRD/rFO87Kx6f5cMIt41H/j+G03Fs
wbpPvZQOoHSwrZZu/C4EhipCazcjOZ0oVymcYk1KJg4NPtKx7NLgp3GWlmv62uMhBihcvJk95YBi
onorx6OUojOxUh/Yt8leYgi/B0MG2CjoK/VLR9DoeiH8aP6bA7M6IeaKBK7md5Az73jhf344A5AH
BSsk37IOdbmXkw+tPhzDOEje9FlvsdWQb5gse+S7N/BCyOqei0F1VlXihcIzptfyL1ExHGX0jJNA
kSUaWfWhgnQAPAAS35KVOolzjFAIZnSo6kZnuPf1aIiE2Uxfo5u2cbA25qHJW7/b604ddwqLxESg
OIw4uIRc5r5BiQhZpGyEKTnjWevqNlcMJPDnH2yum1sJoLftmsLiN+vNtP4w4bf0Fnq+tAr9wEBJ
6thXLjA403fo7l5xpB0tbCyw56ArJjyZcwU6xM4Q0ktgPI/PxO5CWXEtu23onZRh3VpG7TBtClBo
GyLRCX2hdOAeF6YZPwaYVwG8hb4BF78arZFBwCXxxm+51LlIZA+Fphr+QlL43+cN7tn+dMaHuBbc
Y6BV/FqAiO5SezK4nJ7iHIgLPtzA+KLRCFE2wwwMA3KyFD8xk7vTTwGIA2P3Wd+9zDzM/GFdZ5Ha
+9QhH3dODHPfpJxt79TeWxk0r/e3lWwVsbGbH2uOAzNLbThHvfzwy4QZ4LLTGxCGBMdUdymOsREE
768+G+EOnX2AeaLOyit3O+kf4W8skxAPJl8pg729871HKi3syb2X2buQ8CxE4e7NNq3WLnbmFL4d
qh/ig4FWuEcGbPSpzMu/pDfQbyQwMT4JFmoV+8tb1pyPyOp8c79i5SYZiZ8rhZEwp6ezX04I7JaY
7WKo30rsf9/Ri8OlvvKbcrpd72S+D6Xck2JIuKUI7vmXntTZ3RN1P2jPyklrq3icf4Vysx4mzg+t
2NTI1C1CzloFnzNQtZ9GVx8C2z/8K7FrCbFBWToWFBB8kpofhVYoho055V0L2KHIYdQIHtmdScFz
+TsxZjmc3a8xnmSQnKTnKhiDRKyGzBzO30Weh+rPfxULIMVgUA0p2tsP3RpDUR9XDIAP3cUDUsAW
pgVomrzxfAk+tF7JrnGorpaqk/l+0U+pMOp4YI22adiBKxpgCJgdG3dA2HWdRonYsmgp9klJiFRx
e1vuKlL6XFGIL79bQm4mkCP2CZSTGYOMMONer+8rS86HQ2MZxfHZdEBXI0AguATGZ9/ONuM9oGka
J/88lW+Tv+sBKyY8IGxFcUhm0EhPocvjiz+2CbxLOwjvldbsolT9Efy5hjBXqZWxM06pyyUP0yd3
Rc68y1D1HK7shEvWx+UsGgi+HbGpEBPhldsi2fvHR5+ICbdgokcMLSyk+PMZqSWd6wTUjCQq8sms
CmC90YMEb2d7mzwDZ89ZeWR3ZWNacU9RpUAGXplfKS4iKdBiWH8+9rgEi5BPEWy8T4kTA0JU8qww
faPZLkqpw4cdzfpxudFYqIAtTj4WRYrTYPxttDIANmf1vsje8mMn720cPm8S0PtoNmlhrJe+9iiY
mPtV0LC9vO0Tt3v0hWoF1qcxXOznMoWVug1Yc9AkwYjOyeiVgeV4+Ldx60KDUeQhtS9w9IFcFHRA
5J3hVEpfs5SJdOqq6yspLQiAl0MLfPStYWLsMIqsU1iLDjbGqeg5K9i/gG6kE4sf1lqTTlwqQFpe
Nn0WxVT2uTSYUYhRzcyvi/69fex0daJNTBRBupi6w0UNGfCGZBRS2TueEkqpl+92vI+bUdOBaCfm
SQR5uGzP/4OBulFUetcuGLoNxUo4lPZTch0vWhdJB9LGYmc/VGYi5c3hwR2uU6GPCt1rLBzaBwGE
wVlQHhQCprM1bYDPabCcyDKuTljw3l4UxLqMO7C5lDU5WufFHK3CLk9SSyu7/7Z3ur4WIbPA9gKn
1iVGxB33VrkkSwIe7KRRDFOYdCdvPYvkCpMyFEudogiE0FGCDfpXmvS53Hdx54LPSt6qcn8pvW0R
KyjpNq92Ddo9DyDrRbucoDc3uxStacu/D3Rv5nJ8GUFhevTgpE/ySYYLG5iJtlPPWVwg59N6PaLP
kpPLygZbdRutUotfh75lMK7spkqP4gp5PtN19koNVZnYAtJcayTLTQ5sbi31rasDPfHtUjOcz59q
eKGUkXmfzAGwG7mKAk07M3bK+TIkV3mr0ifpDZoRQA81uj1YGQ8ahZEuqLkLBGPSCCwlEvPDEl7G
QYIE57zVq4QJ1NCI6tRog1zUExg6E19KZ3Ha/bbor8dfW/D8MiNO/SHWBhNEAz+U7M3cSjhxQ9RI
ws/JGldN1dRuwsh/KdrNGTeSN44NeJ+qZGvnGfuaLqd4jwTiZ/2vF1orSWQbdu/H3rSsI4HRiBWq
LC24w925W8Cbwjr+eacVoprIxi6hX9OnCXfFWZEiTn/NHFRmOYdJQrGVZRHrJfzZwJxQmNVXWfM+
WyaXUarOUzj7y/hMoqQ4bT21XfQ0vxDISzPvoLYxp8LNlmeOyTbkRW4YqMHzATTa33JSNQS7MOHw
7vOteiJtFFawsDf6PGCyFZEHqx37jr0VnICmSl3ye7YRyV76YAJ8Dt/AneXPeDQUqsCbBodiXGlf
BxAtm2JZSLO38gFUg4lhxctjhbyOPWxkXyicw/RBpUV+lMxlNvUWhKZxFLKVWFichgLJWdIA7fOg
OMV/TAP/5fRXedPqzLYK7SsjqwXX+/BzX3EffrNcne0fbie64uaRTG/PNO2AE1Uyndq+Wpkc97Bh
pHjI+4QB6tT1ZYL+9lP19cTNrSE8bA68NDtFRDkLjMCHGrLnivprgwdnD3lC9rnu+gzlZlWyZN+m
vfeV3t3ExJ2ZMheOo2C6aJx5f7G0hnMLSAOJMe7xi2WMwpFkH6N8GsUyTqhIYDJ+XSc5JEaZhBU5
tS8KVNAFrOCz3Iw6riqdGc4K+um9ugZ30XM=
`protect end_protected
