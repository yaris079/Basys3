`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
C5SP1nrb2YcJjBnAQVeCS6DYuRdEzLBOST3/KwBzwy9ejGxF0Seu5obO1tm5xlwDEGY4k0/2K3ly
zhI45L3ARg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ncZY8QjRR2TG0OkUVT9G6ZcliEHVcZ/GdtIxbL/fdGC7a5EgZQl+MxWLNZ2RfDapPCMtIGV09iv7
OI//sgGR8S9iKV1urktHL0Xj3z7/lttkpjZV3r30vMefuti/HePo/zpymCpUxxFmZFV4maRhMWIL
in4A16PFqsK0xxotiow=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MlqDVwxNgGjXnqtdA+MiZspyvhmjmsTwUOOoFkwqNHmdvkCHO1cFEY+eO9JNcZ7hjJL6dGSi37T+
uFSkb8TLFjUghbXgqaHVZZL/XNjHKnw0vCgWTesat/+BTYbXsRN2TkGlEnWA3CXkOb0141QzRYcF
tSbowwYC8a/U/UTc5+KK54wxpcdzOKstQwwBISc4KH2y+MYXCiFC4hO/L+uLy0ySFUUwfp3nSxPW
65jukdju1zaNWjo+n/c9qZtwF/BRKK8piU/XNov+5CEn+CU0adMjmgJIFjAnrprr4pekhM4N25/8
Px3O9j0fc3y41P7ECcQjr0slRsAe53DAEozRwg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
G7dOE/gq/xWLuL/Df/sWDDRYb4lYklQAg0Hyq2EGpX1nAzG2afQtiX99h9j0robvhzgd5YPOX6Ho
TULSb2HgEaIs0YtNOuLTunUqXqKD5wvL86uDMr2zoU/zErSslTPwlFurhwa/llFKeNv0hDoKdnCi
HBQdE/QRU9jYiuDqhqw=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WGfdn4i4DJiuce1MbDLtDDhcPchtYQC/e4thElQp5KFwNHcFBhASwX7qrelQA9rYQNpUxzsbWVMh
xWskFyoouFDPts46PdW7W5M6FkSP0aoo8QKsycowcgV7fK7kBu1IgYtuaJDvLI/R1N9zkcuRpZEf
WqRTT4xUBntzMBNQ8Z20gfrYidgbOWD41IE0m/isrCpOhflo7GAlple/R3Tl71RDKrlq2YBI3198
lQCDUQSL+SsptcivA/8zKYBpvSMWM0u3VTXVqVfJXtXNJY2hzvMyzOdAMTdyQxgyYgDFuaFjtVRf
f/PIIzjwvp+cBlit/W0YqhvY5VUWWoEXY0podw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11712)
`protect data_block
yBfHc99Y3uQbOaViN2+Sd6JiffYPD4HIcrcwI11bJOVmkpbGli8qgMxiMzXG8sHVc0vdbe/6S8n+
rooczmpCDFzrHVEYKL8nJrUdB3/wwA5247GlXV3DkMvRDXZdfmCe777EPz/r1w3/OTheg99JR/OZ
YSqkXHdC12pyPz1dqQ3/ZJHd1AfuRi4w9dZ0TvhvfYytshvE9c49csMT2ats8qIFDFy94JOoO3SP
YdVdAy3Q81VWdFrbEdn2j/yyHaVeumGm/DbB+WQlcbMYzT6fMg4+lwwQdo/fm0TxpLxgdH3ExiGb
4UXQ+4ekIO6504L3m6Ue1N2E1xdHidpP98g/NdyxtaFqK1vXI5QA6GlQI6rtOj0uJRL8furml8zv
2tbNbnPCIkxwwqJdEzIIw/GuvswXNzndrX9L0dReZ3caaC9A4RwHxLJNzoh5hWpCW1/6UekOG6Op
GN0msFA4vFcv6AEfGfSeaMbgUzwZV7qAi3Hr9moHCmdqJJlgz+HOikPUv9l0AlRHFRwhi9p68XjJ
dKPqXr1DFrjBfqWx00AUQdk+IVBacsDjHRdL+RYMcEdz9qPEX4YWsrVOk4Fn7K1szUIcCScP6Fo0
gPLjaduyI4zEqI5tWrMPLWt1PXecrcxhfXfBi74C0aLjKztoNHNQeQB0FqMZnMDIgq9zroN1EFAr
C3jiHSBc3yi5vC7/ijNF0njXoVmwH0qYoQlSbD1aUO2oTsWcWaqk0++WiKVP1E07Cwzj4lGiy1dR
OBePDqVcYgzXrfWIY/jo3yzjos2oI/mN7Hh6/MkiM/QYPaEBpR4ou4gFOo/p1jVFIMZ5PDMPDsdY
F+UwEHM+9cNz1rWylUHDGMSAMJeh2mr/dRpYZyzDt5mxnQ85fxZfEzUiRG+87oYa/6cKWtrNSB02
X+mv38aq7/B7J2RK2Z3Ta+CQzWRFemADz79eixtPULM6QwwVRnMlHaTuvvVnU9yo8QUWsElGHHM7
RSp6qTolmqGSU7VNmmUQeaJF82m1QLTp1ciM4kI/XbC5FCvBRaub/q/j4b1C85hLWFjAarFhsLGB
9Zbk8hdjWJlT0UxRvYUiDLGUXZdeJ+YLbCHrMQCp1eDi0aq5m6NYcV9Dwjsc4DA7dWNtxAqLBGtI
byNzG/KUVJDGwiDa5BenrQOybp4WdZC7C8n1TOWnn4WpNiH+3iSjpF/yufZ4nLc01yeJGIFFkE63
bqafn1iujaanvTlDCuIveZn8OM1mTr1Dk1RmMXgXxGrukpAgxDbtn+rdrOYucOiZCFDW8eJmWASe
/oXXKSlnOb9FTT4vyZMITrjg0Y2kREj1f4LIbFfWsVdDFmZStpcmeXcLvbUX2OojDDQTP5yuXHXT
aW1aSFO4Qjce5YzFI00qU6aDS4eZeTCGyBj6Z3afTxsume5Fi9GgIiU2o2ggQ5IdebdqZR8nccVa
CVDBHhQicDPeWSDGEm9XM9p5siaNrsnmSW3yoP9B656Mx7h1itGIsqSuujyNNXw8Gf+3yDyvdd6Q
T32656Rus3roPJ3ESC/EnvfjVrKeIrwaUSaJUJL3SXYsuQTMsMtpO+Yi1csZ7a36GihhHb+i7rQ0
dh9czza9ScsjbElimxKl3wgkNB+4ENuJl8gvnsgbED1VcavadjlLvZapjQE/AL7/wqH+hVZhsoFI
XpgYedLiF9q9Xaif+rKNysXX/Drk28IDQ7VNLpf/gi6kljP4MHG+4usfaa6o9LQYmOWHWSjywXqB
8oMFoCZNynVLDRK68jl3DHi+qfic97Fs3S8DROrP7NHqq4eM31TWPc0f1er1H6TaPU0YPc7JmdNK
4/lxc/iod+FEhdqTLVnxVmc/Wqie59BwihTEEx6p2kQqhzaLFb+fKitRtWvcEFKSIrl1x64cMv4e
YEU7DoaV6enJDMUMXGXJu8EerShocZXfGiVEuWel6XBDLgjTLUpAV6OesWno/AU2ad+gl89Kqlbp
/xJfcULV0NfkAsQBvLQfHZwPra6LdmttcXtns5JbOtpRmDRuFiviCU5cJG6ch8vYTLOftBezAD2V
LArLCFnMiP0gCxNIvSf/3S35mhqW4OqxkbFifN0S0m+Fdzude837PXpuyKOxisDVYNyyJyXERuRK
cxKqB2K32ZTS8qB7FY8LedNXd5GwLgDuBrN0MpSksEvfvQ1cGetaYT/wbmr/sTgUFY82ayMXF6ME
/274HKkWcDhqd788LZzYGefDm8xEusVnh54ykSxrZ1xZkttFb4Yf3oqtFoQslVkfhoxeMKEoT99b
BYotv6mCwBJRKxtObYQK4W47SsFndOeY4nS79PoYjuUaiPyOzvLW0D3F/l4uyIqZkUNZV0ZTER/L
mZymcEEFfSELtap5rNFQuqJtYnBGfRJemQjMfCKfAWegc/HlTo2o86TwGbYUBeSyVq7Dk42VQ0/j
/VAlwwpWCtQXXV49k98ZL2YmosDlbzXVyM72dHxzizgor1FT4nBI1v9dWcF/SIMFgyuGfIXL6hUG
3AaiNDUFNDzV4cm/KZJGt72nofTVgi5F23bXp/2CGUcSvzRL0jTdhDYr97Z3YpAq/UzQvpR9uD6o
hVcNTJNxIqAyDMh0o3UsBnPnW4SymCTowg0P6yf97pvJdsuhKCGGmDEmpFQCNSr02mNmd4sdblhC
gTM0Izj8TDJhvaaWVMmrbONUF+BvNpCaxFpupYkx+Y+nNW++ZfuEH5oYGEgki8QMLp5cdcFLUUjx
0tw5LWVKrE22mqTNRSDLibmRy8gGb5rHlQVKioBL3/YBOBXBZYIOo0HU366NNyyWlbJ56ho1EE3c
HHMmVWP94DTr18hh6Z01IOUu+pZK1Mu6bHFjBevCdjn5wNvl5ZhUBIOX6ExThYoytf4JHsEwh4QX
8QpeRe5I08CFyc94TovkDS38DhFUKSOS/pHctFaZhGsj1qFKwRR5iD12qoXbfZC3W3jIKDuPFx3Y
kw4N4hICwSsnfry+WbJ5Sc0PIBC+37A7b0i5+WuJ9hvPtVAHAIdFwpoz/J6NFUACwll9MK7kOSYM
LZ1cCMr7SsPO/4d46tG3Y1f0hZKll+D1Kph6jmSeXYLNIcsEW+jwWUNoAs85/+NELjn4CQjhWzYh
GUbDhJbZvxzMfl5ZKAHXp8r/HI7aGU/bGHZfIa2qsycWxjTuK7MgR4fNcdiLpLqzD7Nt91pyGoYR
sGaBKnHl6GplVgaNACG/HsHT8s6cDINYtHEe37k/3vgCXbn7LM2Q2QY1qcyu7iNjdGupqnYcHQTH
2D+5ORF99eNItCW8ZJn6cTmtZYO88zlqWJ9Ot+mrYtMEJnrX9/YgDtosf29Pc36jHSZJwaCwchz9
1bRMwhoB4bDdhCAVNEfxjqc/sixFcA7QbLxat3bEM3qpDzAAwdWfa1LFzHIekS2x7OlHgFtMO44W
hkj6mvEdWF3AyIRpT6jKlteZPw81X3k4/u4cCe+nJHEltfS2O3Rf7hKsUYJCuPNEX4WW52y1+FXl
eeJeHr1bvA9eua+wafo1xNHo/zZIvqLRJDB7q9I3rSUYZgUAabehPVAtWkmxRmDnWqqrHuvMMQ2x
IG8CHB30087R1jMpEiIerug55ZGUTbIpBfpk1oCudDWpwA6u3OPIv0xr+EAXTQFRoUbTVUQ2aIgl
sg06IuXX6y5E+fDoGG8llujoeeDQCl47NQpmJhosIxGw6g/hyDv4yhFE1T83KE6jgIFFLb87xpwZ
k4GwvGBGVjjHuVTI2LVqSZkXLxfE9IGGS9BzLMf8XtelXPFlYCXfUTaPxTkZdeTSTa1jXvtQspjO
DePIJR5eH7NBHPxr4p4Xvh37l2SecMzzrAsyTnXz6/ldjnWQNv2z+qSaJS6cmMegulkAJpGe4lHN
h5JLA/WSOz1XYgPl0QJD87C3mCMjrtYKaLAIq4QfUknLFPVBvrqrHa+hdN4wDiRtVQ99yRg5nnTW
uDfIIzooV8mnaj/uVETKei6H3eyc1gIjLvzJwIA8rHLWSov8FYvFMqNmboSPMcyvpIsHIzP21QzM
jF8Pdm+mahXJ1qjxdQw3A7lXD55zSjjxY5FFR3IWyS4vPHSx3Oaf5oWssLn78Hey24c6uq7ZcJVV
X0xAnNN8o+WTGb9FGhY6btUtuDGH/Td+eZD/MkG/R6fzHCtDpMzm31zMwUpGmTTOdEVcAtquwVM8
MqQ6sdTQyWMm9sqQBlXCU8uxjcqT8HdmsqtfYfjb3iG2yM6GfrzwX58lD8eNXj+2gDBLEWhk0rPy
IZbTozAbCFQ31nKSJYMR2Ergg8YjohplmGjo+Mq4lcFISte9dCI1Agh1UEXTtDZfBhmdv1sLsotA
8rWF/WknJeRKDTgT4Wdgh63I36LTx0kwQ8rGF6VOQfV27YvfsubFDo3X6x1lNqxAzAoe7lhnLVJn
qOIo49sF50iXuKx+KIxPmK2s7b7iFt/qfU4r80X4wQtsuT3WoQ9U+x6xD0BPzEPsf7LUIdtHs2hi
tnlsPsEMtHqt2r83qCOk7vwgGKexhS/nkFgBz3Sem6PmhZw5HxleDAtVo0KoXLiOJdN17p/go+bC
nud6WvMjzuhG2hatrn4CX9eI+S0nfjARg3YyBanyvc6mFii1Aky7+vLQKn7Jo1r3rIX7JOpszAK6
tmQ0yWC50B7aRr43/vcyl12i+xbO2Z/9kuILM202cnXxBWJRw6Yshz9i5b/rMWVd4EHNRGAS/yRb
pdR1CRkdI7/yWf4OktOQQpuX2vjAmjZZ2rl8CFvCM1FqnytNwB9Dlmt3HAKS9FTqgtV2PCSPY4Lj
7JTk1qRaCyvUkjdGeT/r2+HaY/240C8ooUPYy6nf9l9pan0mgzyEow+Rwpwg7ugSZkGGVnk4y6o+
o82oLkxnpDQOFFYyb4rVfIxC7k3ZFU0gA452snxcr3tyLZVdPcw/OWeK1blQlYBO8xMJP7drrpmV
C3c5crN73yLsJXnu26h7utcEn4Bi2gRRcFwGmRX+FAK+Sde0XWboQP4+cslv9rzLRaRJTCI//YB8
ZmLP20yh/hvLZ91OE9VnKdY9wCOKx9ZkqfhoGSH3lx6b7ZwFYqAuY0DjQsrlzHFfVOeTuBcxkXuX
u/AIv/z5NAHFb0URsD77G/Scl+MS34JFdAFaQ39XBs9uSWjDbKNrYUT5Ea+rsVRlGbaNZCsMH5HX
gQARx+BiVP6FkXTK25CjUnmP5fcRo+FJbUXg9dcckF2LDkkFrzjb62NJi5H95a5WIfGaXUCV7+3l
ycPZOhkv0MRYfp00riOPhT1lGeIF7q1HlURLCHqOYdNQkPJIrRuO1E+qQ8nZekDSTjWzKrkaEpnG
+PbAU1Tr8UOsI0HAOFpL43z/poi85dgTCxWit3CkxbYbRwdWT2smtbEyH0nkXU9g1tjXm78acGhO
b9vDzwFVDR2XhKOAse2rX0h4NEq5TjiKnsGqK0xfwo5/X7J1XvQ7t3nLVKxHKroeXROOyn7hdXCC
0EwIdFYiVb3+tgU6H5aIRTgogCzQLnP2ci0HypMbkDesH2oaUjfJ8XjuWDJdyaQMn1lDlUtgkdhT
NKfSKRZ5kqcB37juVYA2xra3qMq/ktai9fnTFaDgKim1BclofLfR/W53rbqKlIZMUcAWrcSpyn/f
7aNgN87kBMOdP+2Oy7mpa3ghHDZlv8unz+0W0hMf365atrtGf3RV4NfexHQwzO+O8bFfq5HsbQSb
KPal5lFpXcxkE///nZoc7OUipVQo4p+NxvQlfKD4cWejAHSC1/yhofJX10rxGD8NXiLQRRMeeGzW
lw4lChxKklldnEUS4PKkMa2roVwGJQNuzpVNu1pmFZq/84RiDJJBXA92Sopf1hTHvbCG7HRRWyby
c5xc+QbKj/cJ0nRQOW9HZH0UleN61NpuehmFW0iu9qI/lTqo1ukt2VKvfDr48ts2KRifo/h0YD3g
ThwQ0TATvqZB7zYeX7NXt2PMt46x8zQL1XCXZvUArm4X9Y1oLKe/N8hcMNIHMLP9+YxLq+DgGDSJ
TyrPxfKxHNSx04z1phLfIJTI6aO2lyOReBq4eT/+GwjGCQpW1sIILcNCwCf8k+o5Rq75DD/uYui3
aJ/gpXJR8kkYOAmE7n3YzEGNd66Ec+qN+x2TcMoX4fshWr/8yK2jjkP+0FZWp8N1AfqxofgfX0pF
F1h1YKrNROUrQyRcuJA0nH7mFwE1rmmMW5AjXyMT2pGeF0K0ETA8HexVN/5E8LfimdPzy6373aRL
GiXb0ZokjaQ7LT402LCOxBsUd5refBX0oxNyJsHTpeO6OYcZ8tEbjvBdvV57PPL0VfFX+Ks4kIRG
TCWHYIWXR7CXjFl3FiBiInk6djgiaUdfjXGwCeVSwsbJU13BrFN2XvhQXHfB7buaAnc1I4+blwNK
OLVLpjEVa7BH9lCS0FfFmb03Ai6Hc6ZqLihkg26+HUyuT/krdQwXQRnUSieyneXQn3ZzrdZyow6b
SlNJTzy/zzs8yPtV+QDiTOr681FM67fqQ2BHXSkDfOsRuM6jYw6YIGPmPwekZELyH+MvMI5ZLiaE
dubcGgrWPIz1z+CotIOboVpFdV+YjOUkAYEvHaSup2cKFPu574OwW4sR9Pu95XHkHMNuB/okMTwR
u1OtvM3U/mnqDutNJ6jM2ReJYcQeUCwTWpfWLEC3/xbrS4L9X7ivnzobql2aopg5IsZmRyctpdxU
lIS24EsyroqOrcbTCFQTnZqCAwPMYsLHF0MRL1uerO7WuFUTATbAdVS6qd7b2XzukAzTXdEIvLkB
x47dkrxJtyOKOQiIxPnUXsm/wvh5TC+4cETpsHi+Ohp9falBKKWv6NlcFI64omsTG5lY28TcMbzZ
mi5UIa9A6bY3u6QoAqV5u9lKvdQMlv9z+NKuIceqVo6uW4+4SSD85JpnzGEMyV1m9fjtxb6QvQ5F
1VYIQj56migkh5BOw5jXRYVPe69OIrqDzZPp9/MtDhx8IjCDQV4380yJjb2W7xUZCiRwtagUHtHL
yp4O4suIiiyhBpmNxjAsGV8u6+IHznfXScpXnzd42LB2H2dvuwiWjvWWezfDGI5yxtrHPLcdvMsh
bk+m9GNDatFTR+cKdIkMKazGLi6tAZOqL+n1WuucBjo7spKla3a5u945fftOnDiQWZnjGVut23YD
+7Ok0lIvaUEe9y8yI+VoXJclfj7Lqjx62UYZMjMF6lGMzjmvWowR9PYI7ZuAZ+L5VRJD2r0JHtaK
tQMYmXcDbTUDo1cNBRkIQpgB0zkyugnoOcgUtREsAt/60vJprAZGBuAbie5HiBjvS/w+scbdhh02
J5N42x4KbQTsd7jWlPCi3lOAQR3i7ZKWdWG5n6DRVII2nVZerBcSK4S9ObbzBkKetPx81RqIiKXw
lHFJsGSjp/6M6c9vfbMjVVZdrtEhqndk90zgydKVSnujp8uElQRWQxOKB8xP8Im2b1+S8KWOLCGG
gO+xqpti1re9WoBAVSsFdplZwZ6CcZs97RBzx1pSGK+C7QZ7c53X5QulMWf2d8y+uMMUKTWjsUIi
IeqGqEqGR4coAlx3S+gXlldWKnUbcYl0cEtbYEquHNDLysxFC9NzKMt2W8iCVcxkJW56sCXvqxwK
m2MeZ3nvEWmQb/FVczM84r8qDkCwYrvePBKmNdz/VsVtd9cl9RQ5vRmoWZNrn4YomPddpTKTHqBU
waVAItPENfgFmjzX+RdNKj9YSxTKqwZ5y0ml9wA7Qkga+rLDFJwuod4BS5DeAcvhxBav4UaoxFXu
nhJanwl+0YigdmlD02kJWPFWnJBHEwu8FbbGmKP2n/LmB4Qp4/YqiSFa4/ziDvlrvRWij34lfJnY
xCOprUHfJ2LWmONLv+qtGrwSdWtj8G3BNl5sAZmRSL53BlLUlaxCtSqALVlZmFsYLmZny4334nB/
A0QCKjm1srNjdLylcisVLsAPsEd7IHayBVEml9JEg5g3FDonT/TegFcgbPgWCCHjlrIHDVb9RGpS
ZEZrOaNuLVJ7O9lpF3PvM9iQPB1CkYVTx39GnuRGS3EhRT+7iB72lqizFyCPCP9c7Ed4J+CeAVUm
qXSZ52knMutlh4DuWixGWArqnv9oXZNU+Nn+PNv5PVIKDgnK8pdSCWEBENFUOW71n+w4day8pMDr
KZjt3ThJ5kouvy4g9b6Z2bHuLVmiiygEaMgj+g2t2Jm4b1yBbRoWdvgfbRAgWSyaLwzIM4pFLGJ9
EkEMG89EJycArsOM0NZfydyawB86wxVciERjZmpd3awsb3oLUMzeTtINn0iLXCaf6JMse+XlMfpy
O4eBW9WoVdQebKb6RRTNt+gVBeaEfgg7dTZGczIh+WPDDs/3JmlDgg6xr036tUws1sRfnEL/6nr/
7Xor0y4gl1kP9DaKmOt85YzKYqAlKzPUW1alccfR6KApd3/iO3utu2bzs9hQk24Cox5KlpQr1aMS
AGbiTi6nw6Qy1jXywCcQWPKFO+j3YEbouXL6I5aINh1W8pkr8GhixKaxPURjJ73yiBRYPEte4OQ/
KMGB/9RcRQtz+sPZGYhptFXIsSpWwO84AVuHCOD/9YNLqQO2jwlhs232jb9tkfZCqxTyKGY4GmlK
VkuiBo5tzXZbBD3R7zoYnsmEI24NFdVvUX1Pmfyo+ETmDxaami1zDMx1CTQDepJPSzs1IDPuWhP6
JDwhWAX1RJ1nz65RmlhvO+Mkl5lEoD2CCdsBA9Jd1ugWamOItgYbEB/Kl8mnkpspCCpLCJzqvAO1
H/JiITrAr1ga+Q/IUDr+L/Rur9rji7GDykAHh4YXq0OoUIBvXNUtR3MZ20OJva1kKHn/WBxpTgKY
5HEb2rZGSYB31DOyzqzcoaPf87rrUxNaeGq7BVao7/OfNtYhJiiW/WkI98jhJDdhQfCLNdHenQse
DNiUwl3gQWfUJEUmxXg6JdxnBTBnuLjrkl5308oVFuIwmhNy2M7jtObBjv30CpqGV2/PkiUwwXxj
BMrwVA08vM12g7EIUws+5fY5RRB67NQfZqKjJ8WkVPshsvgBTldlPbwlDfLQKwEB1NCts8vy6ibX
sjowWSmxHDz6qMc6A3bNq/AhAvMUPtYBYJaEMe2W9T9517sXgBL/zYYsq0PSTuQqqzEWfspGPW34
d2OWTPo1KKZRpTqv/dvD0S5fN9dCDQtswyAsFA2ObjO132g+1LaeshlISQZR5qNDMariEDRaJKdV
FL8lU76NfwfvFO89EEux3kdkGIGx95vgL5qzCLMp+l8BCB8wyIibPYWbf1+r5JiUi5w29N7rEVE8
WoI6kWHiIb84GbKxpVohjp4k4LuyMyA1cUbXMnFRaEZwNSFvs4FRf5zpiH6PqLZipbqqapVJ7HUH
NYr1ykChRis0QHk2PphI2EeFy969L+UWhIqV66M6hT9adtFe6tOA2Gqh1drX48MFzJkyHSx4yLne
Gf3g9LjeqjHxcDRoNLBJv+n8BLEwM5LF/u2jQIh9wWKU4Fq2iOcxaBYolkIYh7cCpT5HDv24BPzw
4Fheh9K4ZGSylA2dU/FmD+WWd+1j9F6FrmeHjZBvjX5/V+3kDwjvWq7KhHudZf2/UB9nOXeiixk0
uuXP6qmVseI9TmBdT9cebw/kDVbBama+UL4jsNg/0WJpOdjn0kHNdCQHPBv7deqwHFcZmyRObvaJ
WP51W/9oibv1aOt0xwdBw0NnxiDdYl7Gi3z4SCB0c9k/EHpQDuMfVMxe7smClw3EsTE5fzXQU847
Jl3DA4XcgPP+OvQ+3HVcV7kVvusXXPBDj1Lrr4ioBfvKNTsxHCtxuhh20X4MMA2i0u0YbO5K+neo
ik56RizRSyhyKrd1myqmUAiEFYbYmD7MxuHBFhOlqKrNTusxdG60UEkT/jEunQo2HaaE+iwllhtZ
KpKooahmNBX60CybS5Y4KUaiLhuKS2CJJ22UFedHRczLyMdfRpk+fVAFdSDY08CtyXNl2flcq7Ct
pl6mX7iTh4Io0l5rgjM2stUg10MR6N29zDTECARTAQQU1LXb3W2a0J7JNnIIf1vT0Z7TT01uBIlr
XT8GYfMTW2uObxHzfGCV4UQ83tbw1IfCbYMgJxw7q4vagV6Ecy8RseE7a1/H6ZUnEnDcvCo8tk1n
0eqK/QgGDVd8LAOtHii1/DiqbbbsI5tIZl7VJ1TDFQ+qgklyUP8UQ08FamHOG4sTSQmM2EowR+mp
Q8Gv67cyHIRv/e6YA0z3lQg1ZSht+1//MgAlxcNTZBIGJqMX8bQugFnFzZ5ZC4OlniGBYJApgcgR
hBB+PVIw9+okP+UHjydpLlxomdQfVkBpYQgPz9g2M5yfQMj8f44Csi/PXqwc9+dCfCefHKEWjsxn
kMDE2ZRWw264aQe6+r+6iEyqsQAIyXjRQxzQOftrPbHKPjuSWVZTzBnAx+6F3iqBacB3cmvUwx4e
gJHCue5OP0/eG751prLCv4sr4loFwi3uUDvJdrSk6ES9SP5wvSSuECYHNBdRC1Hr65HtwzgzoZQs
WaS2jOD/YSAmsJ3e/to66zmES9HTB337TY6xgTXne8QBSqLM2cOM9fXrKm2wKsB0XOLk4Eoy5RBM
bYAqLcKIarfsLMi1CsmwxyT0c5cuDGj+diXNjldC4OSn+38mMOQV7Np6TqGMwtSLjyJkzwvClEBm
Nk+43ERFPGKF4SPzRxhPFRniwPRpcwgGLhG3ugCVdkE95wMFolhQ6m46hK0syKwOKFTsukh4eCDk
1tflYLZxjPvooX+J5giRmBuhpQfRdV6uBKrg9PTet2Wd04xTco5lWBsKvOydbgTkTOTXZgydCUFp
4DX2cbeVPOpz/xIiFDrXrBcJyc0RXRY6fU4apoOkA8AjExyWyEPB6e5E/bZkPCQkBOCbvPeawt/b
SX79X65YA0FLMGpmbrfxC1RZ4WHYoBQeXBI1bowGUbDkCPlFtC2FWQIZZqvxXTqqrXgSQOVDnXwB
708UFlr5MswDbf9lBv7+phTWAl8FsEeDJrZjr+WpTb/nNtgm4qkCgdHBmDi6e3j8fF63cqAO2X4V
W/0tgPlfGRQG2XKS3YG2vKvX26T0qypDor+Zf9NUFCi2JAIXPyp0+/b+DCeaLEGbqrbdtu0gpDUq
WAGW7hZVSkSo+0uWwBFrOV31tRaLa5we0pVQhxU+s5SoaYimrhv6inm7AIRUlswh8GUcp2J+4/vf
mIClDvFlHAV5KkrDIS5HwZU9rQGfSiRvQ0hsjN0HpXlDeU/yF5MYqS+NMOEUU4s6SVybZvwO9fh9
dD4o8z2ybX75Xc3MO+paK9yrtdA6ZoGuGloxpkaF9wOI2/e7bX4wqC6C3meMQAvE2FSdvXCq0nQP
QR6MwmSfYg46DEew2tdaMjYW0swqcUh9MrEucft0p8P16155XF+Lck71GrpPwaFTG+08NNczoL6P
tmBIV0cJ+rWe/mQdj89rTpObeq8bNvTP3Hi1rwS3uZaIP5W4Em0EblYPjoY8szsBmj5zie0ZQdvj
6Km89HtNiTZtNuKBePGX5lMhwIY+OiNGIi28BQG87a0Sh5x42wK1vT+uFWyAXMkynOvQQT2GBdOG
4qhna/8o1kkjG9iSn6Vlm9NNl/k/SRaJRRmkQpMZK0ZB6T3dZXQKw2TmWiGMkXsvU80SdKpuWK1G
V5VBF7J98ak4Jk0W0tf/aI/AOsfxATKy1Rle7GFSeX7+3FE0VmusTzinOgJW4eaqiUdxZNK/fgj6
5CKjFGrylZKd5/NRnTCkhXZhtHp1WgB/VUXRqXw2r0JbhH2RHfQzKWECBRmcgv/xoWVmFfoWR6fZ
powiU0JVnvrVb16/LfZf2LNPNhBjmLeYcdf0x6U9/H4oau8S0XkMjp3GKmxne9z7330t/06/1ZsA
d9w2NEWQ52rBN0pRcHOF5w7ZWCM56NzlvdZS00RI4t+kUwV3tWx1Baj8Dv0xYcyCTIVAAMF6vjiX
z0OkjBXyn84pY/LFMY4yPkO+Sa2p7zjsBFFqiI27IU09fxJWSGDDXA0xJEcoKrcKvLfO3iC/CcLl
/fh1OlB6nKp6j6x/2uBCcQwsFuy72zsSf1i44zMZvXi7Gfjz4wtUDft67skd6NbcorcSW4cCk3PG
UkSH+bI4uZL72ycjFGX2CddFDUshx8jXX3JmXSP57kQDFFWvL6fgFXXlvGuFUsfoLu4oQQw4jV5F
mB0S7wWAkyOC2G2KqUf0UnMQFzv9JmLMd+xF9cclIa3gwKcU6xe8mjllO1O/KL7F3I7tof7zAyC1
Z3OVP0G0XYXLI8EWahcoYqzSK9uvl9WE1/qW8ZNAwhCtoTOKXQuvDmbgBnIm3AOukdl17GiSQer8
5ZXNQB+ZLCH/GzkT/UMzdU2nx0cHayHzyGrwUkvi6WAJB31IQAcr5oSS5452VpY30ScD4XSOADT/
3HWaH+rJ6wAVIPHsrqdtFoGrr3ZGy2ydMcqKlI4ZBATJXlz2e16MLaGL2j0OOOBxz7NBuQYa17bg
aIyKdGKm6hrzZawYEK1/TZBhoUbKNJoT/9EGqbdBqTlIDfmcyjsK2f3Nx4Ad6Ml48CsssqIDLXxJ
JRFbXHjNjMgdVfg2ytMRkyuLnECh7PBFZuudar/D5YVwOaKHVHToreSxtPUwFyamXTctHg+t8Ybh
G1KCtwU1cq/VULOYn5qRVI6X4rEwGvVDVaIJr+hWFUJNfxYzMIPbqux9SmqIVcoj9nS0ZkBgZJOf
myogSyi99ancpZMLmg/zbKfTJUhj6He1u8z6+EnFsRUnsc2lSSyD2Lka8amZFvZLyT6vGKtDnzsa
gxVLz5/PAcDMF/gqJds1sxnC/nN23pA/sChSLErIpDpEHgu7kJUoxVfPHYXheHh+gyZ93UudYhgE
/5uvagg8J3qKuINg4ExiAfU13ZAUT+azfwakOFG/rbiCFdDdqgiIHeP3hXtJIveO7qTOponGNiOT
+OfDuv7tclvWfMwClMnozKdt+TighiMbGvndlWD/ZGtXX3Oyxo1SCCEmPEFX6T/dC/USMNQvKY7L
1wN0f87w7TpauqSVtuTZ5bkCbbna4Pflyccq93HmPVraLB+I3GowZ8FJQyHas3//G07psvxjPAgq
qrbkje9nNB5I6Z+iwGZQnEvbCSEg462QAd6KZv+aYuztNvmIOaaIR8iTcHufnf4pdn9wbD8zAuVC
HOXjb2vcSj2I87+egQt+4zjbbakG+xHja0MwlKxJVrSpnY4lpR8eiVNVReSM3uV0da/gvTY9ekfI
iyMc4AGSVUlGpEDdC3ze+7AHN5Jp8qG6qe7cCI6zYwmddnw+ZB+wU/elu5BUSy0GUxQfRpIyVbuL
slp0VlhIBxMepTztD1G2J6ODW+9gUz5QSTipjAdGC2dFTxy0r9FNig0v3OMDU7GIHV7H3PoV3Lgi
tgaq64R7Hk53kXlwzRBqFU+cJA3q/676vQWsHRGAE28y+m7msxi6PcBI/VHm4uPioHDRtLabvF2d
rWo7T0kaI56ojYuYs4gHAbUiMPf70Hl+UCrNtBB8aK2AXxDrAsfmjDjaJCwJWDmw8qiDqSxrL405
JRZb0ZQs2jKMLGxhaIeytnvPIlPnOnpB7zzYdGGiz+i1bXC7Z+8KXKzmFUtHEcuZPqB7c96s+kwL
xwTojMm/YE/dxNFcyK2tkLwEAbWl5lzJuT92ZrSMxSxAcbHnO4KJtRQsGwG13NuMPh5EeVn6Y5Hf
705x3HUeWwDz/GHmfg32d3ikQ0ZFoUxTrZb1Qxh65Clm3tDa2rvuqHEQV1Lwi8RnOAPpKo9HP1dg
z3hDtIItR6eBL0+YV2kr5kg/wPqAOzUDgWdj+FQyBWKhmft4gvEj5CQfEngNo+yzBpW56thT5Sya
ymdM6tYapgabnpbigE9Bp4giLTJLx+DqgBp3cQwTW0G7WOpqI2BaZBUEVepJeQaVldfPXebqFZdl
cNSwzMce5td0CZmqHbAJNoRLnuq/kr75IzifTl3fnkrLp/eGqovOPMB2Zp41w2yOpykFbVXNIkSV
QHoCVPUSLlwhTixOHmO4nh04Flm+/nXxOZ3QDM4xZQAqleWpyU3RoFPt6MK+dFegVIf8p2VUTjYW
req7q5ij9i0R5w5YxOIUlWqR7kQH9tc8DwW7xYaAHL/LSkHIrb9wB5ptLsDuMaoGeS2imNQIaZCR
jgPQ3hnnrc42MyXDeY77muC+AgLCmiVWA04e/CmL0/0ijeFqQEITp1gUCd9QPRnvPZlc6WcfpNNn
6e1p7apGWwj6S0ZRNVMOlyzx8Okaygjx+0FMTecfk+lzpi4TPdYahLXXaMHQIfOLpBYKdApajpi/
qKeFBg4iN1evXe4BAPxbtJ5a/XWYySBu0YtsmMa05nlJxq/4AeXgtP8sN4QBJclsigDRMIKhKyVw
BIVbsTqc2nWfxv1ebLvHMBwpLWewJ4JBtyJvsidMma26QPuSjwTzmkIX958rCH3iGZiOmaC/XFTw
Xe/5VxUJdABLhtqfXRdgo3FogeL972fc4pW3QYQa7lpOAE4flHg2KOyyDeeKJHejnNDvMCBD053w
JjV8jdS/NRqfnQMAUiJFL3jOMnfCCsvTvRsDGMvsPb3RVDrhcVTGnzLZABK68Bu/oieQlffqt7dS
JM4hWqu9mMeoLCKk/89rtdkwQarfh2xLfUeandDJxOSNr0wzgbdxGd5vOk5d+2p4IQKtIGM9cFJk
NsbdJkKHzX8Dwj8NICqnCaRF+kTa6705+YmWWR6iyklbOrSRMiYdlpz08NSdLr0SESibE5HbGiVZ
sAqvOD9dEGlFsHq6DEeYaJt8y2shSsU9dDjvnCSEjhoDzpMMkQ/QedXzV5alaWhrJ0Wbcxve672n
PrV3Hy5iZVsDOvrVV8BcIgtjY6+CIaDdHxVBqYxqVp4VcWSP5nNOTBZAb7d2OTvKYAwPjViQ9Veb
7iKyKr/v0ADqlwyCF+ZwLPiwQV9DaVo2IvDGVVGjRhgI1wQSUlpgJNLsRYMiiEvRkP0sKkRRv2mQ
5Uj/M6W3hO6bRmhGKekA2d1UA1q7GBLGTP2sJwiNEQtS0ZsNl6LwT11fzuXEmrURYkCb8GpKQlAU
RXBpMmDn4YjKWgSc/Pwb/uVokdx0xqnBUMtbDo5+d7ylf52c5rq8w3Q5BNfeYOIdzhp7AWQSwjoi
3HKcs9KX24RYcmHL5P8GQsRVHosLWTS7HS4gEoPJ33oIBj5vZAqmiFivehgh7/N0p5lyMD6YIMnk
hHTHFkMUtmoPc/tCGDWVzdMPdDNlZvHdyrJeGbl/gPZ4zlVlTPBkVdwV8Mft5PQrfli0SjuHx9gS
SIoQg6Jd+TUFk2l4u4MCGrEH26qC4TWxyffiJQAdtZMBOpxWtYtfNnutlkbVR2Fj0sSgVYun/HIJ
I4WdfhUjuAI9S6y8nO5rjgcUJYFs3HVI5//wrTDHDHdt7CkX6nYQT+odlR+ps4xHZYNnl9g66AjE
101oithq64q/ZKtgn232x7MhmLr06hqEEZ1y79NezML8Z3/BI8w8DN+qTpEsw6yJtdbCna3SH8tV
6WK2fb1x5MhOkBXqKKrqEdAcoH+jtUE1PKJ4O/qHFaqXqQSHjHpsL46/dXXv9FdWpuztpR/9/N2D
WwvLNAWoclEkz8QnCepKQvPNqNNiqM8qJLAQ
`protect end_protected
