`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ql0LEaQ0tfuQFFwAt7nt4s4gOiwC2R4fB1I74BqSz+tVItjHwaCCVsQpzcnQfE0E7Rs7elXgcHvJ
mcAGbZMUqg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CPAPTGKiWpPf1KvU/IhXL65uQZqsQ47pwQfOmWQKwxCYRTzljQ6LsCasFopb165iT0EIPzNta//S
+72LA7+75EIwj7OjAel7kYqf2P+yZduG3xKpLrs624LuHz/5OZwbX5YFK4GU0bbiJ2EiSRfKrz2z
N57iwhXIrukmcbd+9hc=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J9cACC+C4EF9KdA7VrMyoJ8301ZLa+k07ftpeoAKzRt29UuuNGsoTVp/+fEBiawpitgubQSImv+R
PgTqUTbfaoWA63ZuzrvsRA7JO3hS5naHPOKbDNGI4xWX/YHoMfcEmeKxprqzHtM5KYtwUjGKUbQY
M0jjiz90mfMi2YZ+KuUN2rx0YhMf0gcIBi8yYnoTUiEF4TFuzt+sdJiPNrdv1FkeyevkLZ+Ul2x7
+fOVpUAuEbElVLnaHCWASmmAPpXLO866D3t0fq41sPjQlCAbQ39OUMw7x3yixtUu9WniuGLvlqgY
kojMVQ6MhnPo124slRErc+xi89b29hlo4qk+Fg==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PM7iS8+nL1lgKCLbwvEyb+mHU7D3u42K5W8Yi5rJkz4QsxrIPysaePsQqg1hS8rc82+Rd58fYR3C
FErE0hUEUtCmzjrEUPkGHkYf5TF6+C5Z6uiTAGNHtJmpS5mNh0JQvx/3FIAwXG9pjG3WgFKXJ61f
i6BHBB6itDQyFMqfQno=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GBda/49VW3kOU6BEe7kvhJeCblNgfUcvkKFiJIxs4Gc4MpOK6IVC7trQmAjK+aASXeKo86+uY5kv
Q68QUtTRULvsyJaZ9/E0NhEwrECNSGVQCrt4BpI7f8dT6DP6em1m7bMpYo3oKRnLkP0Q5+gtiK4b
ftqKVhKgL/0zG1Yh+8pZpizG80jrU+/N4NjZ4Apj0alQmlBP91LPVoI0qZPILc5hmyZ9wfch8R6X
8ra7DEWmP4Df0QqmCTkFiZHLXD0GBOxnLzWG3b5b718zPAxxFZeXpH2V91iOBIRj3EVfJ4oogSgu
99k/bNZbg1jqGgCpp+Y4QzY/x6H8hog0y5YfPA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6864)
`protect data_block
XINwDwzAisIZcheUFqVYc2bBCrOX4NEGpUTG0FXv9FuuKbCbNlp5OzU7k/uIVxIp6yq1c7R2KNfV
acdO9ksBUjI+4tDqF+f3wuOFCTauH4VWNOB8R4wq/s3UPLwRGjSqtPCKLEzfxuKxmCh+1mSvQvZI
/lPKKusfNkUvI0jehDpm67witG/NpRn6Y2I0PO81HnqtjN8TtOIjaxittDNekg3a8su9tPJpedCf
Hi/VarodEoklRpx5M4t0rkqEiOVIeuOeNlKjJC1q79zMDwt73PX5C8IQOwWYqyuJSa0R8VpKHZKV
MV8FKPA+LP5m+RyfbalWZXO8Q+ZvGKgTIL/yFN2NvLGAgcOFM9o75Jg8x5n9l1u8YGnJKxJCpWxN
lyku0KzWkZDPxbcL3EJn7ZsXc/NpTtwbZh86L7dqh2UMSG9IENQgPMmbaGV4PKghUoNQX7RgGY6e
AFqo8AIlT/Fp/9yFeh3AO/3b57Dc8qTzkCLGekGDwLNqOubILqCpoVBzp3qJEgwB+w90zLfElzXI
rbkqVPq+lnQD+PljN7819JoK/+t9111v+OoDqHzsVkfRoUH+ruPezo9O8lz5Am3uxglLj7PEIyEO
Wlx1NcDxe2Rl8/fEHz21fHd5SnI8lRdjf0gmPPdp9u9h6TE6TtOxvJTwhUSG8BOf+EsHIU7KVKrE
eSZGBO7Hm1V7gZLTFxYkkFaVWX+Dd5mIObWs3UG1KTn1tDMGINsu/vJLdy9kvMixDyEZX2yfGB4d
4L9nwHEs+/psFpg/a4Fkhg5jUETFXr3D+MJPEbJd0750DqAM0HZG2kjtxUTWAgzRlZ/uKI0eLZvF
Z19KIirrdQrGdV86tM1kzhjIVuPlQKcH6Mi5XddQDc3FKPpKTcIQqrP3hbzwEuqN/UCzcjvtwpBq
G7Oe9HUktZqrsM2VRvnYuXLYMCwPrjjCLQeIG1wXBdfbYj/XA1f1COahJna5NIgDpsPax+Mh2jqC
Y+f2BuFm9JvtqeL/CkrvVo9dQc+8p9epFoaxk4dvxltSjbK6QhDhrwdqj/QM28TxorvQbo2sMuSv
g5XcSpYCMWUhHo9GNdRP+Vv2+MQwzS8gvCp+zL+40qKtMVYJSL0Nm4II7rLpn9iDBU2ecRSQcuth
nYZ1SkWQUETC2hpIha274QmenGib1q9Tf6CZl+91VsWjHiK7lhLhEBIkF52GgS5yVq5yAB7x3JsR
4ABAPPHb/Ly0ZwTgrEf1to09/M2EC5vo+AP76QhdJhH+ekWXdkOrDxEqrqwx7Cu/JLHBxUHBv0Bv
mjlsNOW1Rk4EjDyQJkuMdtxgUTg4aBu7+21i2QfvdMAZ8XVjFuMMK1NOg+Nj69iOf2dBzqyM7hgI
+kHULe6MT1Dr0fYSAVVdJyNj8b555UU4EeIqhMoVAM8Avp6eCyLEI1FDuDXvQLq4HsWXLqVeMcTh
n06hyE33EMDDtSaf/51ok5Jt2vNF/tcPeM8QFK9Z9Pde0I776JGG4gYGH5hYz8nyDR+0o6eZq7HX
iubRv6dT1QyTuJAHGDze1Vi4sctmzB4iusC5219j2HyDdh+h2dTFas5eTUpFPOvoyBoo1phj5SNm
z9VNfsJcKB9EkxriXCM9onfN1+a0oFjzIaz4KG/tQxL5rqIXNhfs3pA9MiHp0wlObJssj+MkLymv
WmFu8E15tBFVwC+Tamq15BbwdaiVnMwA1ZhralY5dVXIQTkyPnrDarwv7WcxaOnN3quVYpfvU6A1
EyFJLZFOVfjM8/yjBfQ2Dq9SIGOvJ1lVpkOW4Ml1I3veOnFO8L3Bt/UPkOtvhiO3cm8o/p8MBUla
5pdUeJEkLun445kd4Fq91sGA83vANHFYENiN/izIR32xx4KfGWHQ6KBwAcZF6jHHjERZnNt6nNsi
/Q5/dEipyiichr+n+GlkCSnlxp09QJ63z2QUfynQchpEo2l14Ybrd6f0G6lp/WNLCZ3RqNMFK18k
o6An6R8Hn0KyXs0L55UjT8m4CKV0jH/hRrCF8idD1bM9gy1MRyorxWobd+KzR2subzboVK87Vu4d
qJIHEoHFAU4PQUNuYufWVQPBLRXW/m9Zm+5AqaVGKAn1CY8pXv+9YV3IAI7W3Q26lbm6kFayFV8p
foNPYylui6RHUoWgmnosmhL1bxxCiHSXyWwJo8OUXb1Y8YKslvJdcb01zp6g63fDhVtLMkNvelBB
JryT5nz7jK8lYpTcrNSL2jy5NfJlVpVoNtQyOfq5CNMmD/0y2NvmaGsIKYJseV5NtQYaa/WDvCaF
zDiNIhGiBLkXXX5hzbvS3y9FM4XqxrT1f8n1FyzyfMj03Ei/b5UTvijfg0wkpO1XjlzY6UnH6syx
F6kexdmvSJTpouEzoz8UD/LkVAdl7hFmHu2/8z+Y/l6o0ve8FhS6xnMcKL2TJsu+Q5rJQIwO1jJI
ZsXFlFsQYDC30mjgofF3FO7QTSf4KYj0F/tlMVjzCfCXGjhqFWBdVom940DudR/+3KGwCbxuiz32
+1HwvGj9yR56mWmaGgxQLLUviiBH3kDH1mqPPWBfOu0+eU0+vL3npKXGF6eU8E4/TP8xQW1OI+KQ
F/IWeF0vNth5WzKekWyCwxWtcB8y3K0dWGGwy5z6XHeR8BR8Aj5F86ajLlgXS4aszMtfdEWNOmTZ
bsCdd2uC8WcLW4PYcpMkPa03thqCNlJz0plxg3pfJsqS+C4yDK6eLiJ9b+N2rBpz6ALR7FTTbx1S
1mkwXMO0AyhzO3GgdfZ/G1clBxrFKqNuE3xBfRDLdvH5EHruvgn7BmU8gpytLcGEkur5PFLOI/Hn
3IspV+jQCNnfWXNcEMJB4UhlnIFtCzSjyy3HWo/tI92pZTWKdG/WKH2EDQcZsa6bSSGtZETzaHiv
oZZIWzmNIZ+uKymcV/3pnO4TGQM1D9OAbKGQKKGQYwF8XTXM1C+w8n/1wWdK66AILDZD1rexbeIe
Tip9tcdWX/yMlrsy6zr9c6Fdfmz/Xnj9K1iTD23ePqYoDTf5vjunMVkw8E6U/qNyJOIBR1mZr19u
zvedITyIKkDpvpo2gTtjD1bFTQXaYXQgG0xAQad5+iMPQLrAaNCotqdFVTetCXcL5weBfGKnm1CR
3tjhJ5HtkWtFJ4Ah65EjVCp2dbfmGNKUlIdW1W2FSqIt1JrlF5oFzxPGSoD0vifzbtdA1npRSQJc
md9YeQyULulLYFsdB/4gNtywpIC5Mu6R97EvqY+3bRxHlvBV4utscOS0bwOwBFhlSVpT4NHgXgu5
zOsygi4IxwM2KfamIPjW52cd+5kkgV/kCN+8MBFFppGisBqoxkOXncE6c5alLFRX5EityxTZL2Q6
kVkKMdxxAJ2q5J+clmwtJTEI+V2RFMS0SXjaciamj7aifLfbqqkJVN3gv7Mf3kH1GBchZqyVke+N
UYMujZztZc0tGJe9VNvtoqfyGhERZ+oco9QTh7bZlHv2za0yKqJEv8pi3imL47aZz5Gyb4oObpbr
HuBfo3fEcXv9l9BVXcxLXsATiIvj8xzAGV9hBxVIY/rW1hVjCXmRj6OWYl0sRgpm70knCDEw6Ps+
VxiXFhdOc0rxw3NN8cQZOH+U1H5GB/6HPMO6m1IEuvBRcIl5rf00fkKdP21cW2Odn9CCSmMt76fZ
dJJ/aUx3pQn74+TCemELRMR0hzTYTZ3zZvdclhQbAszU8Lda1w4o7yn0m5+7aDQ76eSRC0+G9fVu
GwW47rSP7Rdt9ABw7HKO3Sq662XEyEhRdAv3di8NeTuhOlzgTG5HV0dwwovLciYu23uQeDmT656/
o9f7UHJw/ePRQoW2vyD5raxSoQE5nmyom+oH68XcRCFurY3R0s0lV3zqreZoOtb0ON9aWup0ACVQ
w7dFdKrm2DsAtNc+LAda9vXYa/gINsfhiBrRb8JjzhyHMAqk4zNrcEqmfom/bAEiCycWOUQp44/D
eDvC/abZ5wt7jUMFD4oTmN3aMbWeKHIp515GUE6i2+FPzcLug9p0IsgyxOixqkmdnOiJlbcZsI9H
DPs5c41of1XreOfoVtNHnaUhjHr6+8qXPFDAqcBMiMVhJDkfZhwsOqUpv7iAWe4ROGkInfL2Ym7f
Z/G3qYeFI13sU21ZTI58eMkK0bcdWfa1cynir/9oX8IbZHKkPDxCgTb+nNu7n1Ae4RtGmcvAgahX
uNk9BzXphDmBKpW/GtjJIF887e9XWlJjyGUpeJOvEdxC3e93/lbZCiTCDt67BBTNdj0iFekJKxGj
LcYulQsQu10j660FAC556Yr1chpNPXaF2TOZfV0b9bveYKl/JrQGX0bN+7MFeCz4Slc1Htse0q1p
lwfz68f/3FMlfjMuzZZX8J4+dAyCS90BwQMAagpW0jhXPnoPslYWq4ciGXIBX/stFUYVLRyr5K1K
Q+DipVfYGHfp82jQ+acslZ9gixn0psLEDDslRB2OAxVQpsPYR6xXoLBB03yEoYaUiyWlMENvtxco
hfdRg3YUxm8eO7tr1DSlwmIO0aAKpHGdGXF0E7OjTlJiOp+n6OgsKYHA3EKyabbaO0AyXLdFBurT
DB88/N8iYbbQmWv74uHsFRwCUCdGyoqSZ6Bh/tDQXkDEGRd5a3fME9wgDAQMq60f/qFugCPkZr5m
XYO/5CgCZ1+tsCX5l65H4BmsK7E1Ok1AP+4HjROeRCFiSWete1bptVtccrFq5oBIPlrNK2rkjG3T
l8PrLhRUL4IQSqtT23n2XLRcU5d3/cO54cOTsAHpjlGr8iVemEnqRA39EfNWwJvXbeqbnnEitRLm
eJXAy4GPAIRcgVGKxjRYfIa0YRB+KQv55A1XmA69vxhSQyM0eJIWgdJfBnJL3fS/o5hl/SRtlljG
N2oPuP7eNotrmgatyuwoiNq3TCCzk8m5upbTlbZv/uvcYMgwSJbel8rlMltmB4wl4oNNq6sV/bQM
nZv5UyxydrzoZwgdsr45OrW2aJO+uCqW6ynMWw9o0a6aW4nMc9//Xg6/8pVWs9rqJ/HH6oVvxZ66
Q4ieM6OtETAv4oTPGa6qcKOu5lVZYodfai8EktHDLj51E4dspYQveCya/0mJHZG1jaJYhKPVRPzl
mMT+f2u2ctGNUXkG1dh6Ztua+PPiBXg/wUfDJom/blh+9mMQ3lxCmybTaU53TguBkzm2dJLX9xMX
TNCauev59gy3x5APlXvjV56M45URPFuF7V+Qg3AeBGjMNL+fOvApBY7GBugc/xj2660pk0qyUxsU
6jx6yaKfdWrzWgvjbvrTyoZvi5nPkBS9EYfD2ver1wskQj5EHUQvu4Akb05cFRpl3AJ6k8H9qk6b
7tcG3ewqE3Wq3/gN+X1hnk7eIEglNUp5s6Ysl6ng9+pKQmw56fdkrMcSB1iczCskCyDZGysvuiG3
0cL5K3rLY0aVRLBirRH0qxRxoqY/GSuKtTHAAUH2fz5jsBF6GvlVkuX+ePSq9yt/R4wE6SK1nw3h
/Kc7clM2MhSlWMFsWzGOsaUYTEK1GjwfK9WeKMlsG62itRtqF3NmPk77IeHoITKdiAVbiOWNetwV
mibbMjtVCbvq48bliiGxGdOlhI+o+N61AJcWGpzCX/fVep/I6s7b9nLKYI6eIbjWd9MLPUyqm48s
e4sC8Tn8vWSd1H4X1LrweXJ1BWXTSpP+d9OsirKy3FvbZiQc25qCK6OcQQd/7InClrsvJY/c3ShD
HYTljfbu9j7JPR0TtsWDUwv/qvAwYXJqNwBgDaH+RtX5TscQyURjEUQTIEpmf6UwAocWOBhhClSd
IkxiwuWdLt034xXIHmWH6YECZBR+1P/cS8skMsxZbVBB8EQTemWlp//Zh2n82ZwkgS970WbVF13/
pG0AiGff1J+Gmf6TJS+vKJtkJ/L1jAbGNi02H2S4r9Q6pKiNT/EGx/3r37v5CQZoVcSjoL3tkJBT
my+14qSrzpp50JgcsXjJr/QvfdnMgg1RCmDsSIhrtUFd9kwbcrvpSwNLsbu7Xp157DzcDLmkChXE
I1cNntt4zoCX3rL74uXq/pefmP507COqkP1IEramb209RTizgFJNnJh7JKKs0yWD/wa4xAGKSuVA
+5orUNmjaybYNkXCIm5xx7E14rFjTrGxjE0Nyah0jCJbedzEFuGZUf197DGiBLral2EVIylYP5VP
3KfDIhKlQYKe7Y9TljImdCTOgyNxgtgTf66mSs7lRHsWXjf08zmEU/BlSzSDllqhfD4GAbzaPq9B
4mepXA2X+PulQik25M4xLMabMlt76wI0Lr7hUm6p7rVN/LChfdqvdz6u1p/kb0FDGuZv6KnijaFe
Y+bsElJDrvlTbtZWE+vdz//ZWsU5uOKf42cXaOU1axfGZAdKRbviQEAPHFtuXcpdvFkrJ1FFSYl/
7LDb0EMNjzjctw0zQs8AFuha/FxZ90Wtse50aSIM/QDScFLHq9xPhR0q41BdCtJTVs/7QuYganDI
+o0AuHLf+PdK/NRMB/lea6aLtGHfzMaK2K+MVpeW1mZpYcvaK1spasmujVrE86dgbJVHeYqTzjQc
+bOeynGPw+oBAb594LaKHchdqqZ6FAkbjGKjPXSvl7LzK7/Zgd1as7yMfNpGRJvpbB1NRNRtuASq
FsXS07eU1Dq6S4DJOdUyTG1QK1aNR2VsoATuMFTkhVt9cE/1dUphy0NkiUxa3FMBEuZ2d75aBdPF
5Zjg7S5M+n57Q9+19D6kmmjTgRQ7HyT6CFK67A5h5pGsVCsZrNaQZgJaCViA1DjWzGqL98LCLCzv
8jf5G/P2BwW1Q4ghRRX16j/jfVJDrh2JpNjqZJOhKaa/+IJWBX+j0lsEsr3J24yHFAswaOTkKYHq
DHD1/e4PK1mQeXQ0RE4+jUc/CSNNdTzGjNrocXnD2nJxxU5M6QJ9TM7S2LZz1Ye97G8nvrG4/yWD
pl7ZWX1SKPj6jcFq7uKwYLvWgkYVBL6Tt7Uf+OcJJHrNfY4JYdiaZo8JcDm8qOtf1aNIq7E5QStr
PAvGxT7FQ1cHICnN7QG541usRShZrbWzGEikZKPT0mnD4kGY/BW9iqpS/5lr6cdgPyfpJmnvyxGx
smo0cAdxx6xLwv/97tfa4p5w8QVr8k1WowQ5hm+Se6LABqLXIbKOxkyy56GEduuNrQrqCSqNOjhE
pObj0rwZ1o1e1REeV+llsC3qLgPz/E31QOs5PRCc7zetjeGK60Qat5i3mutjDGyc3HTseGgIxiC2
KAE+w1zcbruqISJ1GZu/zopZsDQ8OGX/m+Z7p2Zhyi4BB5+7tDxcFbY0VvR1LNZ1gzaEensT6ho3
255ftfCo3TThLFyLo14GvQGwjaCRxENlPZLF5LJtQ0/Z3MEwgV/FrvsNHnUcDff/+zDQl5/DUL0v
0LqqO7XGq5c2fLKt2BQ2bihE3VRvsb936CWpXO7jQGEYrXPEtCOb3EQJbjvt//TGUBv/+ouecTQH
hG/7JWgpXRqV6JzpoVglgjF9RLymUI0v8PoGxyxt2MgGx+f4UbU0gfHezj8GUSQYD3IVsZAV4fQa
cq2JyUpLHx1bgC+dU5sZb38Ea5yx6f3MZlD0p8JFE48jMQf8LBHZHYpKVI4Ihvl+claP61QdxdKC
2LrbO8Shvt8jdqBtADVc0FfsEFFs6DUufiDMJtlBSv5sfYyQMnLbWQFqJzlgmMyocMcCEVhjaVvP
3L0zWEMzXGXtCZhq4H1TtlQcl2Ffd+CXOOFjtr3QYjBuJIJvkiaP0jetJUJghbihh9reXh679dS2
adGpG8ZY5+U+HAR5XPo/Z2D114Tn2fbM+HayynamTLCuQGNOkIhTb3NI8+v9lY3pCO1YVPJ0aAYv
Jf2GzX4TgdsTQirYhL1IocZF7iPfnLhwGJARI7yLIPNqKqQpZ1wjfgCe9X4U4rIs9vGJUcYovxfk
VdsP1mrgE3ckD+37kRil1NNyAI0tqh3TBOo3zIRL3SnOx2ZpfNTW1R6pAfoh+jJk1zUyUdGIhX+7
HIngxHNhQZ2B/0Z3jSoOR1AeqPm44D7tTYSCGj1FRilWK37z/tqRSbjTTNpxxA8aRcBVOw5CZ2vb
bJhZcOMyzdVlOX+irjQncGgDveZOmjcOEitKSfhIQKFCqmeybFhAUcdvYxrEpGrDJ5U39ZcemNra
myDsF7QCHJEUTIMKdTb3STA/n8n8eqotssHiSQTm/p44kA610c1d4cx0itpUzH0rfW9w/KZJgpLn
Jxezjl3+Nppu1JbzMIie8te403cggla/CcZr2rpPdVKjDI9dqxB1F+Bxnp8GEYf/cX1p3CyVcdf+
0HMkq4vAE87/LTAMDr9MtKozL5kHNQqIUg2aZWxuRL4mB+5rAHOvVlo2zDx7NiXlec4ZNLYFSTTT
mEXv5Qw47QbI3Vo1TEO+gybe0cj42iwg42ILuWZFV73GtWC3ZA6c0ulUM2g71Lmyt+vnMP9XGwSU
q4XOFn3c2JxaA6JGXOhrNocz7cQAxzvJtsYAFa98z2MhqRlYQjSe0L93NA2jdK138IDJMiGC7I/r
A/jkWcuOnh3/ZiFCikTnkKpyQscWPhXp9cjKSKk5HtzPTZc1n5bEqXycrnp6vUPeIvwqxgNELHtU
qbDVeVDnLut/vuC7drc59jJ2SG82vkD6EoFYE+Kzi2EQE4ApJLRvGOwzyX/epHWnObXVh82yBAwC
zskyFQzG0IBmSMDHZDLoyY6syh+63csAEPG5uCi8Uel6pOHwZ0cVzDBq6G+hsrWzZ4FRgT1bRhs0
p6faSjarcE+fr6OIAhG/QmNW8dOvpD0JfuOgz6D7hnh14hkGPi7mvimRybGMGLyymgyKkQ67hK5D
xQ8VdEYbTaXLUbIj8yVi/o3atCLYQ6fFMW0tZE3cStaJTCz6RysZQs4VdMH4J9eLA89zTle8Tuoa
AAzYZaX9KCg4sqMTFooHN70SVKriBZJSlNVF8Pj0ZL0YNwZniMMD0kqE5WYvdSzUvy55TEpddQW2
onjeZyLFKbNUc57pPyd1uydmeyNopoYjiAgxa1U8ekQFQtu5uwGuGXMkX2YryZR45kDnlCM4Z+CA
J/74N7RhRhikTkxZDHaRX90s/3UrXX5HAu4/CbkRVtk2M3snu/XP+hC17+3sLf3Gg1FrJadMyAbl
kk7JrGZWaiE1hmQu6UdzEph2ToJXKUZG
`protect end_protected
