`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
T5kTzWcCVsu7qtbl6i5jC5m1VhgHh9sukLXbgMkRWU4NRZfZAyLu7wLMOK6GXAEX/zADHeezxEGL
Ig7hV+5/Tg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Bs2WJx5/cByzQQ3HMJzTgojSqiVApkShnpjz+86N8OEvKglvTPVOcKDZqSdGtlY/ilKoyxqZG9gv
2ps7Znz3LWB2aQICrmQpyAQlVH6wz3WYjircObzs8f5RGS7/dr97lzp0Yt6e79uvQLiyZxaDKoL3
z6C8J8GwJfgqbzYafL4=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GS69kHkR3u4bEyuNI3HfKE1LeqqDofvbWi32NqA9XPCxMdPZLwPhpDEo5+4CyTVx/WfW6EkgbWVJ
gWKiknqISCkfjsTcuvnTAD9kCad329d+SOSGY/UBSKy27OcMnxc2Roai4lOHpvewV1en++pepPVi
a4jBV9nvadHsHCP/vj7wTZhx+1p2oa4BSPlhZULqIQx+Wdq4olcHy/Oh2qoXYKrE1MogK+9Ifp72
SbqJwpV6kG3U1HCqp3mrMmaBho1hBmjjOouMwO8SpjafiBWJNxgPOziBZYWYUL3Kk+VeEq1qjd8B
axu0VxryNS/xV4sNjZRvyPWOyh8V6iGlRDuc+Q==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vQb4BJ0g19XsYO94/e7tiOkZCVtG/0aLYO70QLfZahmEeM4fyRsFrtdhiXHNuRxlvBDES0NSl1OF
2zf8VSohYQUVkA9CaLXhVf/tsSkThrf1i4jjbYNHTLn411hiEFm56kvf+2zgpWFX8pxvuXlPdk8c
pBRJ4TXEqWtLJ2moKfc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UUj+Rl7K7E1r/+nWk71dHqxgHeWrzFiv/mqnt2DieGnRYecOdJ2aJK2VTFbL6i609rcJ5H1xEsWx
x47RhLrWXOCzm+Iq/3ZtxmsccPMTTXo3GfAxQEYSH5yrBpF2tnmClcuKa0bIKhFGJf+NnWsEyhXR
RT9FArop057D5FtEufCew5aNF8PaK/oMicKChzt63qjjCh7zC1iUXJyqjimOvROqqTtuGVbaVW2B
WCmIqelE95ZRH7i3nRnF+UkGxS+WTnRWMuek5fEeP3xpo64NzaooJFSGI67El5aT8GVTqyW/dq9l
wxQwrbzg0xYbxKDSqwTd5KydpbYU+bNlOOTCsg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5232)
`protect data_block
3pcspUjKYEmgnuibfLAqRldIldkR1Vf6xUqaI5fmOWJuwLyPkdWZ9+epW+t4RvudtqeSlIBqqQP1
D07jHpFVTIzHc8c1J119evfTfXgUa6wCDjTRGg2Dwk0ig5foFyaM1XqdH4ZA+ApFV6GMwonLEDci
NxUlau6xGkV56xkDHrvY7o0c58DAM2kbRQgnHGvnQp5r6GJgaIaNdmpfCIzjfD7mjDj578k9QhRE
C6fHcb7kccNzZJzMJUZiz1BeXvGqugk9TE1JEeFicZX2MNi/3My/gsaPuFrQfenVeI7yWlQNfnlg
TryZdDAwVIzleSPio6rO0xlmLQ7iphXWNoS+kHslXIiC598BQEzohN0PkBSZ4El2juctBEnx5298
n9EphlfbsDTkEdrO4fotO0e9d9v39jjpS4W0MgXQibmEC+iCbYhvOKnUPqj7yX7muJLdC7CQWD/A
yxP0QMVSj6RXyBAEUSCmQLeDaGUFQQs23Wqh2DoE7K1B5A/dtMxAUmoo18AHYO6dGt3atgtSs/RZ
6vKOWCWDiZYyN0erKwcBwNRqpzoX3KX2NGrww73AfuI71JHtmJJOlZ7RvoVf9oQ8vKvHIaa03C/B
wjwj2M4S0vqbK/wuxWdqs71bHfRdTgEYl57lQOkUsYXWsY8NBc7kMelOYaI/GP0MIU7TdHIzAxKi
54dyjO8w283KhDWMq970OBfX1xsPIoQr3u6Z2cfN0F/cRE0PN0oOaCMv56bIehJEWsk8ksQnJTLx
N8CjPJpkxSHpAS6EjNguS54iq/i8xZ0kg8ci0dsRBeGRHhDU2VnZpq6cdSxS0ZMdDHJ9A2eYDG0w
N4OuM/PwxvnOFRvG9Rf935tCUzXLAfYw1Zj1VmAB+EjrQhOceoZJVJRwfg/LktDMKU2hjsKL0eQQ
I1mRnsR6y5oT3D1xweVXxMvUP+397z6pYbCrMBR1dTW9QN8p/C0EoP4B5fXnGt3j2VV53xE4pfEa
zi8+35N6BGybeCCyHyJGwezCaUvSgGJZxViTou42hEqWLZkjN3DelZdvGW4/fsHpEEAw1BGLgGci
EqOiL8z9oky48LN5dP5U0j+u8cHKNChd6L+e+f5dwRp8vR3tCin8+3FCLzmocU+KmKopR1NZrtGB
wAqN6c44+b4VbbL5l1FbF3rZcCmg8qiTMboWYBlZ2x+RX6gJGa9Ob9WCBLdMVJSH6lkDo3mxSaSL
a3gj2IPfVgKcEdEwgnoNq4uUKpA4lHQbMLWY/ueDLAPtfRpoZasWRJpR3Fr48qB/ZUoWIak6kMdM
8IuoAHzQZqJhG9yKiMy6KCFniMbWNP32a8yUiYCjXXhOmZfGUKGNpwle1gB8q/ZBXMzbhJWtMWUt
dwgZw8AdOS27yj+rm5quv4Dxo879+X4QHrRM7OxCkOP97I+MUjEaNfT/Hk7p5B+CRA2BJ8fGRTfK
t9XYSkbdNDtSFqKzQpuEvKLtd75oCoOD9+CmyUEjTrOkX3R0Xvj1QJBUaVRztjq/MYwWGjhbs6wr
isJlJ/IlA2lPxl1HknFxMr37Ncw5pU0GU7nA0q3+iIg7o6Cg43fUujG8oqZx634tM9H3Io8uhrBT
3YsRXzyYsLKfxpCKM9OeRAxfpsJxfdFmXXvcqW8Yaq8LzRtksaaRRTtETsmzm8p7USN3tBuG4dA6
4VOULjR0FE0Paz/8eqBCzIlGruDM/5wOcxtdCFGaWin/BUeIR/ZSG12cbW95/pi/bSygx2VzaepE
Tm56CCnfDYBoGCIYQTPkuuIjsK5FcLNgN1xO3ksg4PJyq9v8hIl9wq1KV00OeDBtKlIF4CoAzIVD
AynB5nsbVg6pxE5bdCBvKAjl9OA0Z723DeOQ136kHGErF5BZkeCKtZLN+ocVayrHFPV92REkXy8z
GHgpNTuDfsnKfFHhM58UFtuYAANrulO5YElSsiwfJDz+GBCfg2EwBxPI0MGE3bapK8PfYy0HSirR
wwQNXv/fE9yQ3TfnlrSim6+USb8F5nBeYcNqfj45/fB7A26SgLpysjUg3l+U7lkhL4FYLCANF0JK
KTnmpOy1m9oGCCV5k0oBG/4isp9lY0+D+G/bWDGFKrJbpA7p6iSYZYNCc/UhZyxMnymm5r7J1hW8
oe6bUIDLffQdVpoOS71q3Fkb3eCzcpf1b4A1II6fQZSOi9kxej8EKi4aDLN8AAXKK7JZac3yiIPm
mtN8r6ZKO72Kef8pk4N1Q3nN7wNMo2IrIXW7t4l2MXfPq72xO5tiC1QP7Bj02GbyMasm9siU8kPU
7Q4Vc9vChr/bzkTXQu3kffwo39Eyk/qickjkVJg7Q6ie1sPiUWmo9ah5cSiDk+vRfOplbItguAmr
8edsOE1/J55KqQpNAlFJVRTQYw9sLJoRW3PtyultfKhlsS8d+DAtaNu+dC7t3eE0svD5JQJYY48M
OpV2jRGVPT8aGGpdxSFPz53YPT2G2LzhJxX85dBVVYa4soo8Yp7FyPxj1KDBYSnqhLuKRAxg1FuF
g6zKvPTbN6N82watmOYrbI/lCvDrPl5UEaGUiQCdpPECuemBYXAGi8xJ/bNoCzKYr/hSTYA+Bzb1
2mJV4U3t5j1+A47DW41c+n1gf3q+xwR5NchENKEz/RpBf4InEMiAnk1gKSElX1L7SL/iaiTXhg6G
kVKwYe7BHnfzCqskXab2iYFVdEbo6IDJtyzqmsiE90vTWSrjeWHeq/qsSfjNUpdkZ07VNF+uNIED
O++5KhlIwtSBq5d6glXgM0FUUll1zihXumlt0ABiG2Hq7p1Xp+pRdolFj1lzqPIP7FrI/RbkXsmJ
FxjG7SsobLdsYLwt5wM+7mEwDppwa/hs+Jhb0XWU9Qh2rcXK8tqpivTGJKtTNKCSd0oxA0btwtzw
/hVKBykezEQekHKBP7RE36hUtSO+0mN87jlm1de1FlnH1yVn5lnT0IkER3PBim/JfxMwfnZd5DBU
x/x5LmNSC8qFUwg7hsu5pkB82FCcEdfPKTZR9JI9YeOlRfR5KiJdOpuw6ootxiuxoPIcNTw2pC8L
nZEqx7RZW9+LaPEiQD24F2rLplOQIPA0vo1XmHPLS7z3tBcC66CAmk9czEM1GerLxudYf4H6dJoD
QSRWIgzIoWMAuusAhJyR1xXY/OsqOf1eey3hPlvxVLAcvYIwkmUl/klceR4we0rug9kcguiAeZ5C
hDtJLG1NYyjo5IGdcee4zUX0iMETtrZ6qs4fi1lPUU+sI1RrT5vgFauShoPQtw+WvKy1IND6t1YI
2W+fy9HxcBfSyz4JGCMKgP3q3zd44zhFvlNByH8vKTewWR2py1M3zUrOA11Yq5LCOIArfJIc0H0y
GFbuxwjqPavh/ytiTy5rK+KjUOhWk3Gi0jptO/031DXhwKWm5/9Y5kMYd+HaGzCooxTCVSUDY1Rw
QKnahK1+2Qua1kVZdSDznUFL8th+J/6w2vwU9i3hSh2Vfi5J545ca80xCUNy3Ap/xjJPc57NGysF
mrvGJPOn/Q2I2ekqOhiNfqphHcD7w1qyuNI1+EwKVUTs1TdwIXe6dQpKbF1Q1/TXBC3kTCIXzb56
zRFOJO/YxgyfEu2JY79vXpvO3E4w897rJeoznUY6kBSbNjQmWc0qO+pAwkPf6hCp1c9CPw+MyUpc
GLDONhsGtx36fpGU0H2vWGO+3BCkZlKQjZTOXftHRk3QEqX8EpY6NhDgAOgAw82/3wupc/tRda5W
A929a8YO9hAx0J4DBZGE2L+pB5xW2ogFYWuExQzrPTB0hgzo6N4kcetWkelZVPvKPPdM5rCkKpBP
LIhcSFzOMO7I+/SeXfmBnF15NcqSo/DRgKry11VQE5TB6lZJgC4jYF7LcWmje8RUS8UfurOt4Vms
WSHuUtDY8FnCH0XcsFuWbAsTEFhvBFbMeA4OYgptLzhPgRsPnhJQHlXa4nnwUg+zNi/SwTkAVnmQ
nllnymSyCuPJiNWdJSCSfla3nxlphZwomng/yoaVE8D4es09mHh8Q1OncvG1vUzCLGUpkChENbzW
9aFszleW7GapAbdIaIgTvPM12elMzv2xa5ctPpZ6WacYIKmu3uZJjpCvtNStq49ce1HPgDHTRtPn
KV3bUIxFgVOanwbVeZs6mP2P4D8Mlj2XCuyB9esPf5qADaz7URD37ZCWnzIIEGqZHu+nsgdjYZ2j
pbxyEkyibRnKuW6pAsRFXEeMvNSHPpJuuwWS6RQIJibZBEbm2Nz1loE3wbwxSSkKaXE8WXJJe3ja
+ZDUiL7Cncv3cUz3vWWlF2sGMIga2SV1tZxPNxVy8E+aKlB8U+bdGI6GKs7qDs1fSaJhzITzCJNh
dQ07k5r8vSYt2nfxkCgG+4lsZNCujhoxtOmGybP59Bgfhusj7Re4zbxYqq+1f8iPi/DCMeSQgQPK
HsMFX1+5YA4wc/7gtW+07TSq9r75y8lAXqr1Z4ghVEM4vhLtvh5tNFtCicuPpT07rgAP3yQI/pCS
HKoaOBoCqI8Wg3zcSu1hFK5Y90AKtIrcdTAekm8hbv8KVhBittGqn7T36ImjNqNGpJQWYxksTmpg
Zoi51TfP/cJt/+pyZo4rpvI8oqCAgk8qiERpMZ/jjAt7cYbQ2RNa8+MGy+vY49rcIQYC+RjSdtue
ryvz7G630cUwkGxi4gO/a4euran/yLUIEPtizBcIC64/cJPSmUxPsFOpso8ebXt5XtCjQH55FKZA
8gD3xmNUs5eXnxb7s3HJD3+9Mv5WIkhOi7mqSnRpsSCyM83sBfD2mvtBIWzephx32gCF1cHuQQoq
GP0ZjmmE6B8rWFujTPYLrC85kepRXZf3U8DLrUuMAasVUi9X9jbnVtRM6KPFksn4SJ4pxo0UKF6n
W6Ko8l0yy+jhzN8qujQm1A03j9Y3EA54ZtQCKhBfak+KAE0ynrJdBj/Z3Y6BgryAPng98QApnuNg
mBkAo4hfArOL4VlObhxfwLhzKstn5HRVurrMq/FMWBDSDJ3KCgFQwmKVnsi7MrbDHGHhY9esK0mr
fWgXmJCsQ7OKbhOZJP9qhiwmEkGtR1ehKKPJzJ/Y+ePZlN3IhT8dycW1o9FSL5+tUioj1r94+w68
bGlugilIGWqO2CRx9CtpS4SHNQ7lTE8ZWwcX0wEqhwgqORaPRKtju8cawHf9oAHd7Gyz89RKqqT0
nUyIfSM1x+NLbMJf/AYF1hi9E8vSC4FUZq27MVDiL7AFAqJILPL5zKtv4pnpyN88pKd9MRZMq8Jn
AG46elGRXn2kEiY1JF76SrmWPGQ2owEzxVfIq4RPey0dGQXeubLJQtm310Az3EoxNHRk73BhLe5V
QB5r1GZuK2AEWYJ0tsLIgi+H13QYQ+4vNod/ONN4Sgvxc3Qf7ZvXemmCHZohUXOmemLwuWOkTD70
UhhMzbaWiRuBawmAKU8Asf1X7l2YFjoIBHKnKNIhnFbuo5TdeNrcXxqEUSHHRRhsE8Y3C+va0h8w
h491SeCctPYRwoap/Eq5zK1h/XEf3LdP7lrU17iMmXMogquP0YLtD9dgi4MCBTikuami6LVYZWxo
31BEqDytN3KLOdRdaCGXPt1PNpXq/3XtOfXnDIWB+YY5AzQ3WiqQDxDwzoUTyuVbgMzv6rNaCQu2
3/N0lm4Os4awbIgH2VgXNbCeV+zRpcXOOv6R5eeqKgx3GFtho11yi7VuVbQpK7i92p/oHQagwju8
LArkQY72CF0LAntavMbsgx7haEg6TlOFVAX28uUAw5cV3u05WRqG6pCLCAfsdVTOZblCjQtwvLtX
8lM5FhKMiVSPOYJq+86qIWyCx+3mhq1idCidA9uimhZ/7K8MF8WSwGvLINv97TyY6hiQY36ib9/x
D2EWpIgfvffxX8amKUAHHEHw6InZhVcl/dXB4sl5G8XOPHieW9DvCLf39TM4zhOwXn5QbO9X4WUJ
skuYtwfVqL45Uhqwluf7R7QLIz6zMQvV0sASNfhSz96qQQpMLArRDE29Jj48vUO99nk+IpN0++oZ
EnQVvPyyTuXUpqauZcJQEwBTIfCvApaFO2yufQ94O4TzfAyygFTd5XL4gDUodJFi3nWOrAXwQsJx
I5eQEOoXg6Jjjq/j3ZLbVIVMVut+5Dl58anOjEnPjGdZl1yu9M5xTmDcFO6lI13DnprhfGvCE2Tk
0K866kacWTQUpIcvTcKj1rmFdEzKwsacKai7tkR275QCpQsOBbyybt/bNHguuksBJnSfAxXI0eNY
yJY/PtZidmdjF19vfHzoRFw/oXn6cJLh0KLRVQeKl4N0sD6iuzwhApZeHIAbHuzzFVWfZV/4f8Xb
HCBS2MQgD8B+onZuEAUvt3/6nLXft1rjo7XHlL/1R7mGzPTpHLIUG/z2zBWWGsl6vvPEa6Mcak7l
GgEdNX5hAHQSqvp6a+M9BSPZOsmCO3opQCPPik0R5+FOYSngiUH17sim71/Y1ku+TLbdXGJ05rPJ
9TAWU8jXfvwY/apGyCq6OgkvR41GwBuHZhIHYFDIbAZ8Df+t343+l7GEAau7PlrdYFbcZu5ahWI1
7QAUaIXI4H6hATfTf7vKNPOYCfKhn2S/pEaw5R1xZCrKgUMGDaBZvj4Rm/NLFGddPKalJt+xfhiV
lwargZBzRlQK55g99oHrm+uPU9lZgnSIYJrHnNmmtOx6X1FVRGowZOh3pjgr2fNmWMaJMV4pnPqx
SBtpgo4UidPuW6m8DDSPkFU9QRHJPlnA68wJXzeN2tED7L3uTxusv3vTy8hxxbDWG3CKRWGc3/5H
gGwjngwt6FLez5OHbTO6pwXBfWJCEEKzXcBMrcvjl/W5wZuGDBzH78Bb+HvnnRfvIH/XF7URAVSh
CADEQmqupvXIh4V0niMGmgyZ0AcEwTz/aVDdxNMRjLhaf8cDFJtM6CrB8O9jDWtJCj1U9y4nmnOZ
vr3BgxevxCgf88CFPrb7hlUvoNHu+qwt97pOoXLy9/fwzcU1KO6FSgGG2BON
`protect end_protected
