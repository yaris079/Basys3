`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R/IU8XltAION4wIJnOCnr20SWrxmJa2zjOsDKyt42+X2xXziZ7FQnzisJoWrIWCSEHy6/uf3PkGd
h9zCJc/cAg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
n0DOURK5O0LTSj5ONCLawOYk527dAifwql0BDa/ZkvNi4idmwnjB/yZt/E5VOAaUzI1ORkND9t27
HzOfwNFl4bFFg46J2RyLca8P+LA4QkULmpO8Je1/5gir2a8lCiaw5HdovP/4v9jT6EI9yBBgWVMS
no6m9dFbCTC8Y9q+oP0=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O/I5eCx+hHIpkdZxiyJ1Lg8XlE6ZCrGjwu7EWCmvGucgeqQkSmEeAhrAVwxtnac8NoOxHjtWEOXy
GZeyRtl/+vm7Qa9QwVk5c1HHOrZ65gHpYZXCucmbhNo4w0Dw8E5At+6+rrCu4xQmzGtXBLWj3gB8
yKZZIKJhbT4u0HWcMa2DJPK4TyWVInoyeGKFIX84avnWeFTatXzLj6WyNpsBXQQKNJMnHSq05UsY
So2D5LRHdNNUH3mTkN6RTj8EXJHpA2IGVhpQpWKuA3o0NFZ9As2J234X6DGj8uPwazY9qsPMp/7o
zIVrEswrGAEIurDPDY7rRoyuYYizxkr5n86W5g==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
vDRc3fA9hujOkBmbSDUzPJfSJ0T8InucjzpN/kY4yvoqfzcvl3Dr6ejIoMxGACrnRx3dNclLD6+9
89qg9apRMzYmfZR7mryQ5VfYOUkUj3AoXcmLCIqxGgQotkLxzRTW/jVqV4ZrX4LSmTM/2u8U+whG
v6LoivCnISSWrCAqB0s=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AAzOa5k4TFyPylVGgcyQ0hGLfIQ02xnP0lsbUqMlRcaZ5pjyENY3V8USfo6LXFKXz/tBaFSqEQLl
sEWiTs+lK1yZdKfr41gqG11uVCMXLcgOKCG0saRfTktTMlcaC+ka14ZR76IQqOjh1rXrsm53r723
yLAN/56U+c4u24LECy6sC8xVqpMuh/mJbQONdU13bLNk7/2BiF3ErvjGQ3sOgCIe9FiGIwdX04UT
OSfwH54yJ+w8JCFJv1XWccZRmbHl+5OPuMLilVoLvczqr3S+ebVfYPFIE85xZr8O2hKSnzdw4riu
kfkSSoyOPrJkTljCAfGUf3I/Qq1E4ifT3Z7CUQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20160)
`protect data_block
8REPtuaSi6b8aft/QdkbKr1QBVSL+Jj83efRTmlxSQ/5ImwWGJR5jqWsBDUlJs+yJlZomPJj1u5a
auYo4bvFjEO9sqVIQ0VAXDpI5BkQDOoSAEW12PDxG/zg24eQpMO0LJNR4EOHBb/fWBqIYVXXErBS
Nx2SLaYnoTZuUBXBU2r+3QGIwYby5fjNqX6CSAd2cGW9iLtzDJTYianRP+5GJVPycjd3cQFkiN88
oELEmHLioVepO1ib4Iu+gl1i97UPCoQPkCPn44Ghv7yrUZMKOBplahPOoU/Puv2WOWlvLtcd5ZNs
P9W1SFVnvWMGsfyTZCPvQy0tBpMQbiwclAJQHbtyL+GclFcVnaxbiCL/uxrt5m/bixBEWXe2OXzO
rnzLV8wyexL6v9Hlrm40uutwXq2NP4YXOcnG+gcwCe/8GAjvCqiIBrDzVmR7/hMIphGvhZV/4t5x
+PM8d4OzEKmCpqa515zOgOzkvIjlpj2wnFrG5ToO/QcmO6AkXmYPQV98EKzZzABrRDvFkSquLkxx
1fDIjTplLZhO9ouDOsqfzakVCxJtK1HYmiT+xf1bjyN1pbe45Hhe1+KgtdS+q9h+ocVKI6IeWhuQ
Kr5iNf+88eSwKAT/r0ZjJRo3Pj9iWerIvZYcaXDq7xW2Ze8/b+e56oCm3VdAVRfy5ZFW0Av2Zrx6
yMtT5GUv3bi+nfchSp6Q6OG/vhZIWwlU8mjRWtVwezSa1UTzr+3OS+kCjasEP5jcl9+InElv24zr
ki2cQb/lVVulmrNzhzxXyaUNvky/v0Ppke1FTnJZijDzQVXRoTx2o9sUjclJR+7i/TfBIiWEbAQX
TqeZtbtyCAJjnOh7BSbeWjMmktxZxiMTY9iMuhKbQTiEFUUsUdtSP29vXe5KmoE5JhRSaUZmOyku
ZLywcUmujMeM7HQ1996VP4SArwCWWCT35tEv6zsMqobuuAPA9z2d63hQRQvItTcacNeJpu+Gd6xY
Ml8zLOvbkP4x7tCqMJxA+hMS4rP0fkqyA1mROUSduC9Bd7ONoyg7k/Mg8EGgCgbzTOya1neFnvl1
LQtsgxzTkeJM8dJwnjssGld7kTA6QK0jt3UTzwErj2m2cdsGzRowVQHBsnZGIuZhpx0UUvEeOF6k
t0pHHYzlEX8MI1l7oRosodRncpxhkAExEAPM1m95MTm5TEy7zALKePP3WyqO/S1HzPPD2PEb0bH+
3kcRckqMdk0BoZXOPGG3Uf1XZ7NzZ/d7dBDwcV+Al0RnQLM43tkxZicETPiqH+P2V2WYBnNHXlhX
Qw6G/43yI2VjxOGFDwZtVqTgy7uO7LVWq6M/3pCcir2t6+1PMSPLj76w8WqMjsi8nB4lQp4Z19rm
Y6+ZkCsrzEUxeuPYog2dB805/ZCwGAWEnimGulFuvinqBtq/hQz72LvtK7HlWvTwzr7h5hbuKE8/
ofvj5t9jDWBggaGCDewvPHsdkwebpAETBtVbPCDNOf/pR4yFVjVTrODit0YfKLIHvW0tX1AqLEpO
he7qtkn3dg7VNXB0phFz2xh8xUzh7UuzGwAJCLAQAqZHVlSShWByzV2OD/vWCCScJjX6l3xBO35+
CCqpX93M5d03Sh1rNm992vfQD3lr+WAbBOwZI5K6lIE3XFrTAnLUa4QnKEs9+u6peNFIQA6ES5dR
V71/1uD75yWOvwBtm1Y4eQ+6szMHHX/81zbTJMJc4FCleu59joP/CZGbTFBMrwXb0O9z21Jun1yO
DftXor4lEO7xQGMmmKguzEDz0KG3dmdYWQhXvx3q/l8IDQ6wYNnHSgh+kHHiTtdKC2cnD7FXiBv5
QK97xyVFCMu1wzlOsRbW3BdChGFBqvlaVcHv5vAve/kPUmEAIY0pJoXdrmJEwk+RRYRndVCGwCE/
5baFjkrvxk+UdFNhWdr0sKOmDcREn48pwaqDdly84tWWNFp73goo4ISEuxXOK5hafYHe8rBIg3Pj
fw4QWwt4717kacMH6jSQLwL8NCJ9Oj5vywDgag4m2w8VXZnHsoEZXDFq1z8jAIYpZZUFq7uDrDV3
IHLZuUcFLEhFX2NeoU/e3Vwe2Yw5p2hEA1f2npu+RVqb2B6ne4VvFjUd5vafKI4rLvcz82j3O2eD
iw0Jb79wbWbIzFovwDeC0oq+ACqRWmDWhEtl0qn4KZqMSTdgT4gP1O2ud2yqJ31TTnStYqY2NsHv
LEQDfTl3vAEROqSbxkmjCyvr9jQxlxO07afEWbOLQDg/Ea3X4GdxioYOUfqUTLBRdyNt7gbsW6O7
d9h6uvax/pVeomWPBPrM3om2KEqlrUTs38lvCbKIwUJczmUHC1kSKlTU9qPaUphGklVrY4qNX2Un
/gRKLX19L8Rk1HECXPvAC2xhHNjTOuLmFeVEefa/XLBwPQE2AY3vfrmdxy3Kr+k6/T7l3MxeEh0R
aamlv/iXfCr5pOKPI+msKuALCeWQTZyDiqA0VcKil3NUeUT2o19BZehky3D8ApkST0R+H0d1wZs9
9Bm8oAsnWWbkx4DpqyrQFhWKpGa0/iuukT8rD4OS3iTaa8yDnxxLrtpMdBeIrxTTZP/mflvbwPhE
8qqXwy0klWD1KU+AqCjN3GXuoBdEu5XQ3AibtadPhlNLy1B+AURvwPSUNnxZY0wGfNeOjwVp6/FE
Chq3dgisnFtXikL03GdIPco3W/g6dz9YQMe34d1g6jIVAFGfYSYjjP0IsosbuG8U+bB5sg5wKuC+
SovnOxmSXPrpg2Ev62Sy3NOhdU0remubB3Vkf8KWL3X7FuPL1Pgz7vJgcQM+DH9WzzNZOWAMsnST
I2q0lUeC910I02ZYUjFJIHavv0NKdET1Esm49SgIIIYE0WxrXPYqA6NwPnCUcoWAVhGhVE9/XpyZ
V4ApTXG4KbrJOT42rp8RPSMp8LT8ru6B0Jf6Pccuu389JKBzG33jjqbamrTmQqiBW/dZqJgMPd+9
j9J79jtKGLHARne98lBQKomf+V9B9l/+Qkfziy9gyV2y9vKE4P5DTJSxg/8jBIsJFH6JBLxjwJJl
/G2VUtmkbmWD1UaPlzKYUcAxRhDIW+e2zu741fUyu+aA372xLXt6PHg/gRJEgSAOVIZnaCV/ru+B
/3RHYjwinmXHHYZXq7mrGHXEGmgFQ5omJwDGXRSy0tUnqDC+ofZHAcQ/xpZsqh6bjSr3RQqPMHmg
qP6v5Q5b9nE0HT8PP0A++Dwpv2CIqnAMmKczVCx2Bd/ocajQ+vuUx1EqVV5QYSwHV34bawY99KFv
WMraca3K+9wD2IgelkTgnDOURObM7/lDLyqfyXEu3OeD+/5OICNjENIpf3/sQlHMMqIhJga/3TDx
aqxo8Qwohis0nTnjYBml5f229mEKZ5QSdMDob1UCzlNe0T+IsS9rbXvM76yUrNWF7pQyFFKhG6wI
G4NYOSjUA6TT3GkYB/4JMGd15hQwUMqUFZEGmrgHrZ+Z9zvK4Bpr2LWwK66xJW2yJIGheX9CFsYG
U8NBICsyxvaw1s11IrePu+GpHLI7QlrY8sE0dP9/Jky/3FzFtcGmRf8NKPInSipGKtOVzlZvxyGN
am4/Qin9yrHa/cxME5KApW3+aNSyo5iOiUWob9yhWZeU0xDU6gBeXsX3r04HdoeCVPFlQnpfj3qK
Kh7AISEKhRavd0eubkY+iAHhmO213AvABwBhPCOHy0yfWAMb1aVsFyOObm7107ymVVV5mAFnqBJn
Sx305RV3erumxdhIIT74q7hOmNd1CoBpOWaazZxtP91ia82o7nxBWFUlYAVYxGb95WyYQ+d/zE/w
qUrj5dmknS+QFLX6kNyz0wxzmjBzcFtJseSAezq0Gl1D6K3b+zMDG03rsx2OWv1UI4KL9R4BG3Sc
4MSDcSHT5l5X0Br7UPb+0k2LqDrCscH+9M39xIL5E4khfyAd5ifLYbyITWqShaINH2kQ6xiqnlxM
/5jgiCbx8E9Ef8Kkvmi5g3dxZdTPfUCIUn9hah9LC9pOjI/FZCzcNSdI8p5LYidPa/JIYNlvEo/w
/jNDK/G5uinYpVvscHrvaDIYRJO3zdXeMQXWdI0/s0BfFTroTQeBh5oQsRhvhov0apefuafq78QP
YE2PpibwJXOdqZWXyDj3YdvIqUB7AoxWXFHDmUiuucNPRSBhYTTPUky3ha2vsd5cLVDgRvqWWSdB
bgIV/ppZ6Ilco6kHGiZLEWPiUv96Z8DA8/jJ4xzDHwg2Sfow+Io0lo7cBVADH4OszRo93mMFsxTm
EukRIQ8UGybDCNoLh9mRPHYEHw9zpYZgxG+VmP4u1A07QOS4zhd6aCqmr+qqechHe/Jlsg4S+2fH
4ZufHjTgRk//CBLGs2TEGRwUT6gNXfQYRjIuUdIKMG5Gz8Zr4Ya7HgHsYpoPCwyKLydxycRINdOk
uLCAOB+6nMtDMFkkX9XXsvSiVbohGDAWs0BGh3ncmCjLLOFdG9/Y3sCaaVwf+og/2GlTx2hb0szn
CQC65C1o5zw3cuTa1ypBsQVzaKyJnZC+XuoIL8XdPDap6XxCtE4mDfdvfr24BhOpugh9vViAAWME
4lWAr2dCL2tfDyfe5osd4iPwTs/hwOfrnaVudl7pOZhvHBalATMEvRU08EsnCXJ/ADTzwTNu/Mpk
f5Xgn9EGynWJ5geoiUlty/PdtZLXRcJKZdjzp+7JRvnEWLm6fmlNypf3AGgLCgqQr0XQ32d/wk6Z
ac/ZuH8K/3fv6MvR2OKMWYC/+91dq2yHUqppvqtjfA8/s4icuD3ipM4gbv5pZQfa2c2bnx6NNFq/
v4VxxWQasufkbR7bgw/pD/VrExdBXNpd9OZwkg8t0t/PdteRMvrJyis45JNcBCkZmKWERQYxEV3N
0PuOdEsD/D0WIGvITqWOvYVrp2kQYVaiAzuxJxVdLE6M6ZroytPagnfbrBkrBQugFStGWZFe/2nn
4Lzy9xKfUBfVTGvW015jvZ3C44Ltgc6jxueBA8eNpit0nLVaOWAoYvl3f0S25syEvsLQYw/vXkqG
+lHEZ774TNE0DA72dYqSdfp6lGqKtZuvfHb9nw0I36EOoOvJbRIonfCXZ9A0wF+KHUW7Wex7NXip
8DBRXaSABmEkCGCw8XCX9Vh434URkbXBZxkumshpM32OdYtJcDLcWKOczdi8y/EXgNBGk0KVAwUo
eefzeY3pvqntIDyhpzkinWrYCAc6DadA+t95PzxaXE1ZqbE+rC/RoPYESB4cQlHIDMZ+9YjX0v8I
VJmPPrPXQx9lfVHEOs0XtCePyanbBD+Elrhbx/46k/138CevxsIQ86mx3YMDxSrUPZde6CoqHaY0
3galY58gd7E2jZV4qZBlzHnELvTrfCwSD093EFC2b2bC1puVHYNA27Jjr29DYjqsQSGryFtsslAe
q+TkJ3dZ5yhk6vEIvSC8ZgW9uG0rjbEgahXOKgJWfn/EwalwGrBPb06kNmiKXe5AE4dc4+qXpQEs
YOhA7iFFASkFs4AoycrmXeQbBnAeWGH1+ROGb3tmL6K1hCcOVDsIHE+lM1i5WoMWTjLyHFp4ol8X
sH4stdRpYX4HRxv60v7/LwUX4faqphS4AIufTjNdYIrqCPUSq1sB7yvqQDC9Xl3435B27gWXV5kQ
6olwbFRXJIPEtyQgYltQHg01II1Lxl34p1jyiFiF7jzQOruO6tTcBXmMNC6RIQKLlvAWR0VOu1lL
/+r2yaRUZGEru2261p4MQM98MStkiJrVFIIqK2MdB8dvAVvRUAZOeiJE539K9NwOlWN9pyUqJHZb
Vxrdr/6oyxBGPXplDYMGB2xfMAWRD2qTnoealM0yP6AWHUl4MH1qwsbwtviuKnMKNNuoySAvHpWS
s8oaGhmh7WXRNyMaW4ZmBEZDHB0dLNWRva6LDkAYegt2nCgEDATo47W12oCxotrLlT7QItbozP/O
r6Q9eWX6kPsQ39bwO1zo02QOFSdOM7+SqMcK9NR1/4qoFwE+yXXyfY97YBENpVGVPv7tjbnAQabO
6T7i6wcpkB+90S+NOgUG5AQ2D5gBv6HLWm7k4Xa9qq6ERlRZJ6Y0R/PUHnpA/9ZVkCTGMJFNuwY+
vXGxUt2/lcC2MZX1mNt9NyeSNIKCIB3SMNLdMjI/4vYAKvDxL/5e17DzctIOZvnDkKqs3AXQ7Rgy
Aw9G8kLw2MDeaZylMGAwpNJNGIbnKBZWkUaR6THRPxXXOiRypBn9tELENN5IUuHLomGSWWBzGdYP
oRDcmudvuKdqgpbk5GEqxHgWDTZILicX8W2FodJngULRbDItKcTir0gdcHk/obO3CWU0OuUerrOl
Ju78EfEOZ3bZuPbC3x636db3wxyqXaZnbxqBmJhnw9gLQx5333lJPUGOPcH4gAZhrMBO1tJUiD+t
/kUE1iWfzAxVLzFMXxrL+Vma1RTSyybTpKiszK4U++5NuNro5l0EocYlFtph8p2nWkFmobrG1USI
w/KjJdl8KGu3zXAuYc8ZEtISvF65gY6/eEMgCEMVYxvwAgkrC20dvk+nNS+kyyi/W/56UYd3nsdC
P1TFzUyQogamcOugZqV27AbGhktkJvZ7eN28gxanRkLBSi6FTePL/IYnysFbgsxxoDmQA5f2S52r
ve1wOUO/n+g6+eYzgjlAqW+I+7jAB4Mx8VML+RSQ34kEMjfSo9FwhaO1Uvj9McGT0Q3cEMhlBzPW
dmcZmCPJ9HSSjF7bInDQk6LgYWK4meFAfFYkfjZhx18f5CqE5YiVziqpxKeJ9R4eqbJV6jfUx5ya
WvdAU0in9zBcRcdT7T8KsorL6jEiYnKGet2Ph0HHqg2vY2+WIcx5olrnyXckOArkfC2VfSfDi8ep
Zu07imyUnh5KvvBQ39HloX3MTz5iMpnj73OQKG/puSOf7m7YCemza0bgdd3OJY1hziVmBsHLDxUN
i6a+WXG+LFM7mdhKpaG0VssuiILAedfafnYCrSrlHuEwdrBeArOunmWdDoqS1dClEAklpUduG/sW
njVpfNbwdHmke4LAV2SGGityHx/2KGN2H7HOcpqqA4+Uo3RE7OTAlaD78k1S3sy7HR3SPvaFilmE
r91UoMppXhfwtrH/bHZNPv7K9pK4v3IbFO2kL2qFC1RxvhwIY1ONkYE17crOcq6Sa2hiFpUsOvQ+
TRVxLMxzTLgOKr4jZjhd8Js4J9AYUMZ3l58P1gJgQT33UfRBWiLu99jRPuOlbPEKhyBvYYLBAaiy
zCLF6u4PIshtAqXYIacv+h6hmyrci+RwLGse0b2mfdDYZiTTFcPfEOKGZVVR6dA/XPRjI4/1F1U8
BX5J+vcltAHiMGmRwpuc+rH21kfEbVPTdP5Gn4AdoOAkD1PskWbO4WGU+lM+/zDnejQUGpfql7CH
SqOFbAJUvLhkmtxtaBHwMSsVtWMJKIXZcraiILlLnB3YxcMwwzNNOy/fYtpPRNDC75PTxaZ2c2df
p42S7yfP1xGt6kJ+jkkpanbRvxdxKNWL58mmvzXLKHOer0E3mrMjhCdgX6a90tT93+xBMUssjF6r
xqcZ5att3QDkbcDx2LgFi3Nzjq5scMEI4UEf9pw6GsD7sZdh08fsFK/loVLcqtmS1vLKKAbhlaP2
cU8DZnAc1Tks3ErFO19vPIv2mmlmoKJqW9WMBxHejTlaNwZomLECXLV+2BkTJ70vxBz925Z4UgBS
wbnlPuJXdmquabAMJ5OpvngpkG8uScc9Iy7L5N5cdIJ3houX6+HP7DEVKdgH8IIbgQ5iW1L76oR3
JWoFn+SxphIWmKPVHK4vGhUeGCwB/OSmICJURakZalpPiq1tXS/5LrQZhaYfdyOPeqf2vRXE3x1U
WGd22jvJ0QpfSUgDtRHhKFxGQPVPK08Nw/Ap4aL7/HItVtPFg63xMpmaACQkkuF81MCT8yKrwtIG
nyNx1+ra1kFjYe43cUpuEQ1QvOvCCO6D+ksyTKl45lEZuqQOajqGasjDfSuSACPtFEy/kgbaerm/
hHRnNZ6LtLOtiWNsleIvIjscwUK8jv4isIR/c/WEjTz2uFr9UKNLCorAQSHSTGeWnm2wOQ7zIfUS
xWGWDWIOa/JXPvUYh0zxBg2nm2hRXjgoQPfCJ6cvnpdkQ/lk5coFS/WPvumfQm3DzRvEDfSxNrcx
JlVrTkidmy+dTXiS+f3I8YwZ/76voh9DvOlxQs+gKfZRQg/DYPjWVD9kyZDtPU72Iurxcp+4DPEV
0m//YXYXKeTdLfahS5vccEqm7ahmqYFLSxqvLBx9RiPYbSMuOACsK7Qn9e/DBjqCNoSn1wqxHuQr
uH0mTacpkssATFT0qyzgH55WijOSy/JmsIhXq+q8dOMBikGtWykeaIlWzfzsDi4oAyqONYwjhic0
1sn5E8bhNSYXSnRmtxa2vQ8UVBq5DbPhXGq5q33CFlDfXEk16pQDDs/GdFtAQOqbnzNBb0APmLtc
iFaJkjiF/aGRavrWslkY+7FLZGqhPbkgz04zlPtjXWkA/+CcEhFsXYq73Ec/688VbZHzm5lFw19H
ExcjdRY25+hD7XEppPZo+I1AM3vs0vdC9v+vKD629LhPBJM5IFdA0qaHdsUN7AyYEDsZgJVbEnak
J0WMumZbu5H5IFl/P59JJhmcyJdedfaJhTYuLEniUpmbIo3mamgrotq7lXvMKVHMGwjNNI6V5U9A
09xfgUL2yrZbb/0huoJLZ+t62PjW1W2PRcpF6K+RJCIvyHNirguscSXlEMMuDP7ZKBGVCCrPF0HC
T3MeNmo4XzjdywUeB+4JTW/B0AGj24Q6hXVgaVEjA2gc3+HbCpCPrlV3ycYzqu6gbfoQDoLSesL9
/WVPdZ8qNMTUDY5Q+38P8kZrhkqO6MvxT7hYqByoSbLtayTLGsdetOJZEBS3J1/q5/GJMdhRGJub
YvgMVYawbueYhsq02EWhBw/S2YqPml2LOKPUZ0CzN+H7sNGswW9SuSShuEaTN7XzKX72PHjN9z/T
Xf5byNVMBMtjm9+dOzWKktMrZM9ij3Dl53PArjszcMfUIC2aeOY7jXuqUMN4IwVxq8CIVrZSajLw
ujA3hhowmauxP2yzTI35VQnVdd5FXkE1xCf/IpYplcPAUHDI8mKfcCdMiz9iRlZgMZic18BjB5Gl
9JRWvAI3vQd+m0ROE0tDjDfQhyhlFMgFiGs1KyOM/DcsZksM/apQAMKXYLF+sfQihZtayeTh9z2O
qJ9RYr2tp+hVZnl+LquY4QlWiQ/vV+QOYNQiJ/UZgK5hfHnk0hXqYdOnMJNsXk9Bd5lo/QC6djNj
GAi1c9F+66uTGHn4n1rI77w918Fz+JphfLleLh5bjWD59fGSGyh8uoNBKPdPT4TGPc42XWGuSdYg
vhG+7XzGT7BBK7mWoojhzJquHKPer+3h3cT3AVrd9vXD7wkgaxxGuWt8vLhj7j9hIhikzTvy5WkI
AozKZnDVsUanc8pygZJY+kgXA5jeVBI2kY/elAYYzC3r8YLBowXn01agXnTkGgCuiYTcMU7gf+cV
eikDsWT6nyiP2q0K8sPEUvxmDz4oKXEL0Gh8FSssgEv6Tk3hZkty3w5WWSNpBTVeneLoFQqZQ1TM
OHbTk4HJ7RQ9h90Oy5aXvphXXuo2M1Dg9WAN5ieVU0v9fgcvRbf3JGtSaHnbflptrt1k2QkspX7V
VVUr8AJtFEccs3e2C9mE1s+rKSSDfVnyDZeTj75mABr3vb4qPBM3TejGwSteHsc7b8X+1XlWsQdP
J2mPPFxOkeXVe0+JVW2X/ilv4ad903bDT/SpAcwdRV3xtpQsKmcgqUtVbC8PwBEjika5o2SrvnFk
HqzkIZCPPwnTEGrg6amsu1YMKttR8oicTUm+9FgUqUIhQ6joZkMHL9zDSFmgjBJPQnJT8ahv8EGD
Q0EzoUgSbcvSMIop/9PR+V4g23RXWiOtD4xq68uMIRzZ8rrHOEpM/pdrEMmHgLxn76cuTa5L6u6i
umIKejuX/9VWY+X9crpYa5aFoHHksyXWf8HxEy7iFHDNNomj1HyW9lSTvwW8iOAjhGiA/YgWke7Y
e5w4cm+MoHut9zROBJfNjIcdn4fC7wEPtzysVGZGM5DAsL1ChXlIS1/lzSV4/HcTVlL89+5nxHba
2rBlMiaIT13cj1eP+75tJdD1ShcgJv7kqNlBQJsIjmMbRa5efFNtcC0gxJUOfiZ8LWmX4Ez0Q4F7
R3Cb6zoJIWIrIZf9dWGQxs8Mp4AoLi6Z/fDfIIHHzYwy28Sr4UUd8llqM3apsOcqtwSCveAtb3bB
S8XGBiTC4yyN/iOSe9KP1i7bGtDhCVyOd7MLiupSR/gbtf35a44fdqzQV64hNMuNFHcDbTjCBghV
kOFiUZmkfUTqFQFeeuY+4HqFXGdnu5pEqJlNc7OftwqZTOj6uUUzRBA45nHyTlzV2I+/9/fyX/Ib
CmSgt6btlASIUCtTihJ8UjfWQGTBWo78R9+RmH1F8h4BD/Gyb/Fx8w5tzKiY1zNBBAj8s9sLtBj8
aUA/lJ0DsKpMQYULJlrjeOx1jPGxIkwq/QHf6Rw7xuq+4dmCDUNv+VEpgiUcmH5mhYRoVkdyLCsj
rk5dNr/bqC5MCiN4/KjtNOlOShkHRii/zHjmgl0+fRRvpEaURi+9D3/oJBHXOPIvRnOxWB4wYJHe
+G3jfoKFxrxiGIYKgwVx+NJlWTRg0A01M7XrGW598LU7VjtEv5hXFXo0W5f23F8IgtOfpRWwm5n6
W5LNv14s9JQONcY+3HzqZvIZRu8ED1iemtcp2sDeI2OxKKpHdmrPNQWH6zQrx7OzyQFA6qpgqLaa
mMODyQFvyHsi3x7xtkyzz8Jk4uRUZdk9lYtlp127Vs2o2TDkWW80zTVqPTW2rBsGapVCS2bjgCKq
CDsneu4+sFZZslxFDGFbkleJzP8EW2nR4YjmjLLBMhoJkFY/C1hBR0GMJ92UGe23tRZcjEjjF6I2
ETdQREDZwuqcCnWChnJ9FYoFBFy586yONxp0YoCRaN2sf3hwcQpbf/MclTJ2GemweXduOJU6apto
1CErOenroF2Qo02CKSS6sjCwpE+wJz1kuAj1NJOY19g1gsXp1bLUmkkpB53PPZPe0ksT3EZbRjqF
JLLPU5msI6IRGcw1hH+y9DV7d/Ty6TIl/3cRs+0IOqdquJhIJ6tIhzB6ZYMVCndvGCVewmmEfQYc
6R+5nj9AIliIvzYqWeE7MizXfW+n9aJNQUm0tJQbE2IGVu92Z8OJsBK3AVJXhdwPk7gQ+w5E4etG
bXripjuFB9B8Mt7goDyArTvXS3G6mJNbISjW+oSR9i7c/xJfGNLxGnSwoTwhPiYFRaSOsxwcTs37
jCmM9bBkjqQ96oPecGKykODbtb9HJj/OdXg2JfcvAvZOmomLzSWo0aB3qGT+hn69i4NapECglGn0
FuJ8LdUvSF2gnM6i1ZZeW2HrHEwOUqrz4vf2B96ZAwbr5hqaS/fxTOljB7ClAGl3LnuuhVCOL6zd
lrPWQwYFcIZoNxGqbzVvQvTWgC1gTzKEXLmdzHy5oIuitFIbjCps98zkDD4+gVrjidqVbexZpOX6
2SDg7e21FBM51uQ4Gk9XwEvXctvTt3qPhwIUi5Et06zd8O711ivm2PCVmSzoHtgZpR5FvTq3WkzC
d+iteeXl3UYs0B9FbHnNX2kyZ3bwfhewhdcqhwiTKP/mIv+gBUGBNoEFDu6IuggdMKbdF/piJ+zX
MmtBIlCOMD2y/KHW7xlYR7NW3UV8u96AeEzMhmgJVbD/OFRWXf/9oQZyHT1c0om3fgabtxRI12zK
KQvDGtqkbJ6IQdpfGXp9wtpcYuhzQDj765RWflRDl9LR/ys0xyuRneTrHqUhrvVeYfvopB8/PKhl
cmhVIitmjBZJlIpAd4PkS+c+H+4af+pFVehYfM0LcPDBfC+v+n6ydKPcM6AOYsCeC7bJ6jTQfbwU
V3PbqTs2+5fI+WT0ol8lgYXLtAsF/Muf/dbLypcS/J5S7OuuAuF3HltjynCXQw3+eJ5UOoQSw8Z2
5++apzripFIib0DDkL6cOqxMlYAh+o+6B7boi+7kpwAqP6b7PeMF7Xc9dVs4wU2V9D8CRztGb7hf
7uwnjWp2qrA4r5DSAMeMoHUJg92eMKxOQgfb7Uze23yqJVl0gogUYQghWsObwisBI2Jxl8COuosZ
GPOrDj2cU4Ggdis1NoZqhuJAfjfS5nfA3kLG4TFA7DHSFaFkQ/mYIe6I7nQKEO07T2/DgFvlFjRO
x57IXL25eruW8H7UI1JVXKB59FkH8UxssjNzMyV8lmcVQ0YKV0EHz0VubrlEd9BEpGVP/IJdqjZ2
AzCG8z+g8MxXSvCsVS3qND+jO9BeldAiFMstpy8hLvkGOAoMUiQbPq42zmAzRz1gJhlKusGTLA9t
2BhkRFKbxasW4n9adpyaf3BuBL5ptK5HQWu3wh7KuDPsjlXMxd5ZkWXkV1XTTyJ1eW8psJjB9MnM
JnziWTJe7tA/C14EOL9pzju1z30FGtn5lftAfQrpV3b2J8FtZP2HdqdR5Uih+CiVSdrSpC69qVRt
wo8i+kL0nfXSWowf9Ib88+phYYlKliKyxRBJLey2nYcoR1OAK64EkbLb5JhpvHxK28L3bzT0S5Tq
t2xZUqxxnCRR6m2r/P/4kDL2PW7Rv37Lyrn7+Gcaje6vPzQKo3L3ca7oWYugcYBXjU1xeK9e6/k1
5Ytg6/O3S/XMRJi8QJhgjpFFUZFA+tkx5OrzzCSZmh2D+xkTlkScjUQOYs34RxQXn90Xg8F3gE35
GJpunl38kU4GMlGfyVNE/TuqDUPlIWBvcIhxL3QpY7+7APWpMcOOpnCyeGCdst+luy1Eto3JCEN1
lu+hVO3c5aBME8liloX7BX8OqstDKHAYXxN4V8qcmopGxAzsjTVohHBuSBCH5dcK76mEAObvwYbq
4EfgsyiBU7gRvGImoYfwGgGnFi2PNSsFNnEjDQX+GXUszRjAz9mp4KGOAiY7Dp7M2rJ7+TUaIl9v
haTN+kBEU0edh583+0X2a4TtcDvNsizNDXttmOaXU70dpkzlOGdPP1NO79Se8EqVh2zbc0NBcoxT
zR4mkhEcSc6VFQDXnStmRN/fpk8vBSR9TSSTSaK/0uYBUwu2K9naueRbE0A/xUj5M/Egm5TK7z87
WctiolkVh8cg1Gjk8F4qGXZoe7LWFXbVsiFnnuxVbzWuWdgRKpVtvtbBBDiTX+06/CYUAgwToJhu
dmwUCW5nxB0yYvCGbKq74qi6XQKF6Dugfqchix2haUngFhhDiNQ744RQ1CVk1whwHQm+FBjTuwM3
KvA9+Q8whcIh5NsNzd8sSFrmPbXy6jAdw2uN6RUbADoYxruW1cfNiA1+RGumJP31oTtD6qLM4874
ZeMo1NyzAuAkdVlUs62pYyaTkGe+GJ7/GyXIv/M5uB/MKnGfUnfNZG9OQgcP9y3omw/sNVtL70rk
QLBrPAsgLZAbPUbNCO6waWtlBoaRPH4qBu0xqKEaJcMFVsDq1yxTeG9lsgQ+zBnuN7BK5Cbg8fUW
0MIjd+Sz+1GQTF+zljvJzVGqS9+jT+qgrTQE9hoXJGEFUqtc0Il3LziroiWG/iTHof7X0kvyXhNo
08U7KgIfbI6QYmTNnK7XLPDFikn6qVyQYXInp7QZ3qAPdjWa/Akg6kbDEqvFSJ8aUgwRuwxjmNpR
9EmFW1kxiNyYj4RB9x79AvS+PjxIKXdXHPxW8Tm2qWMvuaTLc9Dtoils7JZA6x2TwxUwAk5CivLM
saBRPNNbe6NFFBlWX/0A7BOvIt/qs4ldrvieUQtUYX7Gg9a60TffusQwI7VY9YsSZIfcicsTlv++
k2Vx0KhfhISCvBUp+uBVBHi4jIzoeC6mrcpTik2FqsAYpVZ3Pp0xqBgN1FNxI4I8ym4x/rQwouRT
TUo+FCX4FXRSFBB8T4kJnSGcpKa2H8tWtYd6Qhqm1lCoU5+NxaD28ei++onH7LeL2zeVPYJ+MmKQ
HFtmJv/RpavCqD6S0ebwDfGjojGTBptibHgjJ5gHTt1s5VnCgJTj3M1A1E1JXTWJ8hux/iy5xANf
c0KBPqLZ/Fil9w1zUnHT9iuDSep5gjPEK09T0h12mSJvjyVqX1jDiMayL5WTc+658234LWlIKkYJ
6uKarnGkTnXHlAnpHjGsTgoIJfaBFZZzdevJibAHFA+yTflLZFgUlTMvrm8oQ+7kHdRaUzVnrTTp
j/ZONHc4q/SFLnatsrHjtIkpdnPmHFWP2vTog4rnJPlQa5ET6nEn34qstysFJF7NcXWs4om5V+tA
Uq58EEDBvxwN2c0ZsekYaDpzn/Z8jgvzt/TMimMcjiqg917hmIfzHMyKbUrgPN1emil2NWtsKmUM
wtRqj96Gi6Y13Y9nRUNn24NhKKImI5NYh4IaqG8Cd0cl/ike7tYxBi3iuxd3CiiyFNk4wLyG5SHD
EmOrEW5Oi2UBVIA+958G0WbDbtBqfuGzDY+xZAPYeXyM0jDmDyI8jErY+aWsWE2zmKdWJjiG1ovU
rF86DvZnzoa8bNdLVglh8h/EcjrNPC3/pialUiDn3XDrM0ayItohQ4sTeTwe4WMtYJ2M4X1XWT/J
/kHh4Op28wa+M5gFrmTnkpNlIZTy+mr3oV62ryuk6nU9BIw1Y0wKgCkMmEIyDlS/eGqbpAVRTwpg
Hk/WGoaIN8vYr6NWnvUmEUMxWy4kkDXxC8PlHCL9WNnZbuWPEOzUCasRCg1pp7xM5mpxdQ3WE1sE
NcKM9KezHM10wj2rtCaWOZya0gYMPi5gcZmQzVpiqUysMus+1tXUBFTRQgAnS3tpEdihVcvQFKpu
LTEvYQ3V7f1zlTvG1lXp49B6WGKAIy5dwsVvM4MWKThKDjetaO5EQthlRAMgOVsoYV1VSWzUWmSA
1FOKs9jH7HArO9BhpbaLwOdPbOKtTIRyodUs7r9eSuABfE/wqojxq/CZDSfPPZersy1odbPxjmTL
Bzab4cldnozxbC5OPr0YljNAGDwrfqdVwN99rAOh4Mz30sWoIfwggDV4cvNXnV72NLATO1kbHqL7
2efjX/nAzSWvWvQVtk6YuluwUmJdfpYrNreiZZbasNoDysgRNGDv7Mc+owNK4+HxGmsniugUDSEW
oj27uwYyjNq9//Me0GOTO+sY6l2ZtOKq8UUGQdu36fjRQpL8CbB9J3dG8QhbRqkujj2oBavaBpKP
RKgUotAWcZXZ5mBwJPqC/OMZly2JgBemvlRtakutxxgTzF7kAx9RyHDTt/DFDK2AD1q7X7Frw5Ga
Ks5Nw/ThlO/lvLLT7iEiB2UGFMyb82y77nbSP4yaV0YEv/BWp4zx49tJrMlvSNPsoEqFnTe18xew
0SjWS0r1IlWJnuE1a2AyYYr9rm8JEIjDBkcV2R1uZiqYkteZuoa8zZdOnF90T/qPvR7I851+4j+b
F8gx2ZwSD09jV77z3K8SUxtwgt4rdc9wUuKNWMa2lQirzMSvIWygvtthRqbUH9MQIWwOa8cR9J4Q
I+JY1YXu5GD5mIAdHKGprb0W6BvgsWbSGJz7yeIuKQGJsP3/qKn4WOPQvxpho9oqjfdkRUbgx9V1
C61WFwzr4rT+91P/fcN4LWCmr/kPJ93YayjFBXsfTKWLsJHCAvkpYtyPrc/os843ETmAbUUl6qpb
TkBqYuvMvNGYqXFO4UBStVa1WrLhlHDK1IcGZLswp0N6EzfyjQ2tuIfT3YOfMJe/Z0oZy4Z4f+n7
5+ByQaDC5y26x1JIlBA2KM7cqUyj0/egy8yRQVwXiyw/D58pmto7kw7deiQpld7ytQbkW4EDX9uG
0euPfO36w1wBbw4ISPDL00z7u0BvB1GmxYSTXeBpRSODYt9kVtSOshHPLZhhKjqJJ1mc/wn2fVqK
NfPtjwj8NG1vcQ2p1gXVES59V3eH5IsySRg3TlbLQNsi7oGw+u8Ox8p59PrO2+gXEOG2FXKUselO
swAKXSe8eAbxOSa1az/HGzHFayMp4/1QbAUWG6hwXtrRlDqFbyDTn4I/S3kxKOwWKveWuo6yHlQ3
jwdGg5KPkdAFdSPbOqVHPOiupY1DM9lr+8kjcdA2lxLk5oIZO5QJ1MnaQ0lm2xGTJ1iBehnWI2Gk
aX4DqBNz9qsxPlSxH4Pkgmcrfnuc47WrbHNPsmzWDxfOr6nefozcLJpupZP/s+w7tT95XGccoC80
rtyME60s/WxNUW5aG4RflkE2VijTDJZxJMuSQBula+H9JUMsSs2zv9bYV7PfmPqiqxU2T028wRVt
kP5WpFZsqaYSLLF+ViCiRSxhH2J5Rf0+kOx5vu86xclV5wJthqsvnrk6NY3Z7McqaUBSEB4w40Gn
rdETjM23CVSGIPOKTVA6vqxR0WxlympnxXilU3+PWihxWImZ5024HIS4/XgxH/F4LME0jGQvVBFw
DTDcOfns1SXToXTyIf9AXHQ1fxSwf+EUwpdiLY9eo/c+oD8lmAr1vt2/Gulrhsk8Nms+/8q7D4W+
BlPzIMi7DjkYbdxijWpw19tipingzVjQP842/8+AQaFAYaiCBxXatcuW4/j1kFW/+Ujcy+WNY0M9
QzoJbh9JXNr3Cwo0TpjLnwN044rAmUZ0zwRbYPB8e3kzmtDdmFBXu85NF8oODYPRu5vmQ5jXuET1
PsgfODtVpqTsfRMvhdGBMltNBACHWa8Ed7IM9J6AOZ4AX3dFtrWvSoKuC9ysVa7GC9spr6hBNJ6Y
7wtI2tvlkuHKPKLAf9TA97Bv37TiqTo0kdrbuAZnBpqbBwGHPUEZJZSmOycPirf8BjpYqaGYnq5i
RiBln6ZzkYq3UBhj85owtiNcshRH8f1GFsrh6SSsbB8tc8haM/WF+IboKCelJLYSFPepJBTJzCRh
vW5QGkLJwwdI7DtNnsEuAPV9jpQJIZH5iTKUZ2N7+pUGCqIeA/LP8SExspKwsEPIlByxk3cyNjjF
udSFR43naK+JO8t07g7WKAuo2PQG84iE4b/ae0iWy2yImlIX/3tkHPUe3cnCpfniieVjcRnOqDsN
vInK+lLx+ifnrhN9Hj3knrp7y573gc2qilNNsDyniMbWaXJv2JZJXVFCbKo++IVyy5IappJq8EnF
xo5n4vuW7fM5DeIXdy8mEa5d782Tuh5SBRTvMe0g8uzAIItsEnTWPwE44H7EWKiPfbC+S4v/Ins0
4Up9LmqOz8ENT+Syy+ssNrmIJSYkv+ftTbW98otbMr1z1FnsBIzJDPWZ37ISaU5LeDv2UfuhzuPO
Y1XIZCtmZtcVs6RChhXnbzRf1/66ZNDUMOooXWdZ1TTeDn2MKpbE9OSX4YTAxSshis+WiNl4l1jP
oa6zqhJTU0hv6QaPks50p7yI+VI4fVs+s+r/edvH1iRhKuKYgLfvjoZUdLlYcH6mNafwFVh2p2MY
Wqy2jubElrwG6YRCJE2Or5QYrLJTe8KfFSV24OcGeaOblXxZxXpFfgsMlCoQ6qQIwBVIqfLyY6br
qtcIN5qK66/VpfzJkNgwQ+gvifvJjM+Kpoco/TsBufVs7eb22abIK+JXUOO0Zg7Tm2Y20R0sfQP2
pKtWW9fTiL++IZIR2ozkj7uWOf3JBMkA8V0RBKFCiZRJ0d949y0sdE8qsvEPDYnvg8bF7Uy0Ag2K
4WnZ/E+Zjl+o6oEbX/8CkgCi2swc+lZrHeFBRDN2MfNwH8uIN7//yn67kdzndpZmoyWNr8L7Uw7V
8LV5oERGz6ZPghCMbFZciXIpZ0o2Lmj+g8svMUvy601VuWs3d6ilaE/liZQHonqvS7I0KcH5i9sP
A5aTLl406NGhFtCYyJTwdF73b9P6wZlOgoZY13THK+FufpmqdfKq+6tTKU1PmO526Wqt1twxmuo9
cyZZur5If77EQh+9pOxe+g/vS0XqzXTnSkIC68fJnpqGDu+htJZFDm0U2w0Ss5DYN7XSwt1JG8/o
XWOUtvWE07fzjhsbcaqVTaxRSke5OWsTPPRJWNhO6haRYScADlOnvY2Xgfc8y2aQRaLVoRqLE7+8
drdAxVVfuxGRuBRTEOXE3YfOoBVynHm1nE39woHWs+oHQkLvHlQot56YKOryQs+2c3SC/xsShZgq
U2qvOUyQb8tnWZ2e/lBxqWse8dDNog4XeUKBRlLEIVRCHsNP7Q+vPr+1mSiJMlfY+5doT3JEtK+k
li0qWdAXDEaAvUbbbw3d07tIO+/8B9P8G2TuNg1sfWfUgqmkzQRhJBlqg2ubqx3KeC4+SALzDnCk
CIKW3PFAIQ22uFnBR9b4cOZfKVmYC3WCJE1f7kFbGgjQEdC9yOHBspCxjQkEeU6U2MVjZgFpwbRv
OqszIYHV7BgNdj6PSdqOgVu0hDyj1cofM0bhDRGgFYyyGbLlfjHMvMB/i1c4IE+RUKiqu7T/t7If
8PSZGaqmG9G6Fa1N8PtD8Ul3yVCc3FblKbGutS+y/J982hdfPgKo3a6Os2vwMkVwT71Y3+tentZr
f1+YWusJbdWtEw6DvTig0rTiPBDQx6UxLmrngi78PhvYONpQ4D7r74pYzGbJ64KEaA2zSr/3h8qU
J3QTxotauZvXgL/XBOpMmieMVTIuvTSnt/P8KHKcKhDdDKMXnLHsx7qXbxdnpeGGr6KGaFoPQIQ9
JccSYnE+IpW3G94KCDV5F5yOceWA+RpdJTrRT6wXhtrvU0K/V9r3IA7nNMiPJNaV2drXYm7ciJ3f
JiQs8BAuOkMHh52xAJyzHPLnhV+JhQkTzkcGLW8nPSNmHi4IXLqgjQQxLRMjBrZh8Yk9+7VxsmoV
QvkWN1xUv6P3rq8ySV0sX2uS/mYJHL0Kgcmq746rdGO6pxgVFTsRT4jYIoM+c0/+DEd24qkpbZlB
3UXrbbud0LqgBSpJ+0/X5Umrbh6QA7znkFkpla4huBBYWuPao2kIWjdd/auy15aBHpmHzrKxJPwD
QDFrJj6JHdq5PTU6KZDVcFjQj0NefaJUFBTxcJLHE0qfB/AMfSiwCf3HZ4qiz0HwlJynQfbIlQtt
hC01/ZIRqKLffWvkJH8wrhEzbyGsPmUhWBEp19cH4byMadYDjrsp2mS+m6lKCTWPKXW/rCAT4xhv
2mEoxEr28sHZqqg+Hu6hVb8IKwqF+uMwkioYgiCz/xk2BxktH18DRrUiSkqWq72VpieExKwVcVbB
Ir5AVtEy6QvmzMklWjiRLy/pASp+owLaikXKD6zfgfIswLQOnyiT9bXQLjAlYu4qFwyrLgYyWDZn
pgGisRCJfu9t2L9TBreRCSCu62j9EuW/Q9Oe3xTbZvl+t+MUIE3MPQH+RpGeLjNxRMmCeb1DlEAm
nPIvyRUPjHQD9n/3BRlaTPQQ4fakqtqqjilfKD9LRilHzQjYw6qPYSD/XTIYh+D4p1GVOKSijeZJ
KtK+WLrXNEKmEAHllI0XkD/sXOy4xdswBrT68nkmbUDxlqw3UThr3uWCZnabGWoj8zAUbsVo/pE+
RAWz6XoXMQ26nmlMPAfkLDhGl4WfJ6SlkUjKSiVLfRYkacZq763VwEfoMFnej+vH7A7DNfjUFmlN
IpYb+K2xi230mksS5tJGDBV5iQd04JQi3JgbCdiJqn60whu+oNUCxzfgN6Gc8XmuLCwFphrvTkOJ
amSndmf+E5q74b5hEIYpc2gLtA9KB/v9GxuSpBsxun/ygvfiXZc/nj5zFnZr3hwQPf/2BcSt1IBg
oZ7gBq9w6e2vTH+JlQeJqzx35CDaNBD7YY05+nXdjjrDynDnmI+RYzs3Fz/UeLdiTur4EnFUHlMZ
UTcHM58k1bNPmv/6VVqLbPGxjQ3EhZqekzFbVlo5huigkL7+O0BtLM2hu94p8To49wOdF3DKZwW2
w0khcl+z1kJ1ZgIe9ZPMpoTmN44iALDitX6fJojgl9FBADuoz4NlnEm/Pal5iAmETBB8cM02EsdG
lSk9Y1N0SJCpk4WgMZic48XzbO6hteDPbiamOPYj/ewuJMF3XWIHO7zTpSTk41JhgpPMpdWdtGCk
8ySkFpOCc7WUK2x4GTwiJXoJ3DHQWK3V/XRhUz3wDWr+JeNsN/4YenEV5V1UjrfhkNhNDcMHLv8v
IqllZCSo02cDy1JhPl4z7Z6cnsl2mI+G5KrFE/BjhikOlP+XyaztwGBNi9VJqZmazdQS2RcsBLmm
sdenVI62Og7OThiPBL8S8TqbsoPuCKVbvX+v2W025ThtZfhHxruvoFOhFxZpfA1L4Im0N2D3sTwz
yXAYyAzYEgnFum0ZrgiHbf1NCeuMFVJhmuW0vNRWDN3rCbqc46DN8HvLDkR+6AlEm7ZSpClcWBtY
IAmJ6FPV42AbhdRXqfmRjIH+qMY/Rs9//KdYhOs+Yzve+ibTfXRbYgXkBCxVMo8WdkO7sOsS7qN6
37dteuQRrZBCIjswJPaXkzH1/fXcXcKyxGgd2uDUEPGu+IUorFPM6aVRptZPRgR9EV2nnGDfjDas
JXFBr6Oc0rvbkGv+IyTGxICMfJzrsZXkXx/NxLHfZ1SBXDdEitmfLh3s1a4rjaFGreMDLoxWj3S8
iAn8TALDkjP/XsbdlDa/R/TA6XK3dCpILgO+CYstCkvvMpa359OnHQCx9UOuVNLF2zFizR0AqkDH
ur03TrENtBgRAboum0iIO4GochxTWgrkiKx+3V3AUWWj47uUgOH+FUfURWMCT3zu0TuDmMtNqb3w
JFPH8Kpw1DhNnWYv8ipf5FcT4iKeb8Xmr9YOVZuXOEpgujid1kdfsdTbr/u+4vxK9QJgrjLu35fh
L7zuxKEZ9IGvLDfkvviD3tQEZoKiXNJR3G455xerVoo3kiE6qqB6B7c/j7RYqz2RMec5+9QlSuK3
tJTu6Kh2DQvqXg46FY7xnml06ZHXYM+zzl4sSqkx9KDQGaeP0/lVrHnvnJjeVtzUSNs3Izv8RRGz
QH/YJJ6J6+5g/JJzAr5IL5SAX9YjFzBxoTV9a9HQP/X6nVuNSYh5gsnk+qnheiiDLSd++xHUDHWR
ZKa9OldV5cOBuXIZbDABHukkfKDbIIbLnsfEtqoJWevCGaGs5jfyXPnT+Od91kyqOgndxxT2yjyw
RxmSqXEEKIF90ChZNj7BLVOUFPzQWZf95H7CDKncxbY5WYIOyLmB8aaZ3EHwXlTiwvzXUy9fhxj0
V38AdK/NPKNiPxfZ41uZX3RWzHHG+kvb3QZ6ab5Tbsd8Z3BCSN/hFe2w0vaeeHLvDZ4FewWpypXx
FziUVcnpMzOD6zliHGrdCDuGaCDZEesdoojqBJBK6OmlmOUFgUp8aGZFM7qnodM6FdXxglldYf/E
O0WUsK5Cfd1JuGFPhyQ5svufSeWvtsLX744WNPMcqMrXcXHBMdFIoN1fscCK0d6wK+E9nCXqHOd8
Kgo/Y0UhP5LV1hvcxrM3excs+76Wnmhk1+TQUK/3DJCerrRaAhBolzUwwUbClR4BnioW/hnTKyXQ
ig5ro5Ysn00WlJocfjkzzV0Upmi79KLIx5UeoXFjnU9hlB47G/fGdMWjstHnk+d6/OUK2lvQvlpQ
NICIdlbMN7JIRgFgWOrt52oU4J0c5gFXysr7OvMpXT3oKlgundPZP26sZ4PEm+35I5PDnNMmbLzZ
VoQiC3PZOKcRYAMg0i5aNRJiPhA4rT7DVe/hCZMk0dIkycpSvG13BV47bPiIbpX3glZmSHMPiVnN
deP3IOJzks6JV+O7IiblHx7/3XeOByjQ67Vi8Jj8waubJaccjo+Z7RXHSas7PA1O9qVLlhG5kFSf
6JVN6mqSdkwKJc+itFyJAK340phdgSEFLBSFQm163bIOcEXaZhOYka/Gw+NaU/fyHQ54dSpPnj57
o3wBP/FkNCp4/GlkzwR7RUjSMgiPUpXu/+HCBt4M8UTeLSFtQX3hJNpyZQ5oC3EO6FcDAF81icKY
j/FEODW6nOFS9FsCkJ6dZhP2ol21IuUEPfn12oqWlL1x3wptrUi2j/brtPFBEp/3LdVD9PiC+U+8
/I48tizSzX/JJjXoAW7SsleTYw5uPYgM5jHoLyEkIf5nKIebAFpRjcchy8NFJaj47WotLgJaJMep
87t5hc5Ele/Cx6Kjd6W9Eujctr4bmqPYAKFO13wA3ge6s05MO164s41ghgSAQxePJS/iNqCe5q1z
Zk4W2oo4FAkqbfNNUScgYLZ9EjxCkRAl7kRx/q0i11l4lHyXXIAB/mxvqc4Xt3/hRuHISU3aVJGK
CzAU9YTpo0xtDxNgMXcP4UWtMG6rfkQ+zULfhLA7edk7sOEHLoMGCWm6vVZHeiml+EnqXVa5/qhV
HxdHo7HbIJH9UC5/SD1v0OetAuEBTrzgs/CZf8FdNtMhuMKtKHeVVsVbxBbbzx8nCjOrjpB9wUXC
ZM8xqNYKTAxxRb4Qy7Em7tVFzNZ+VnyY+74AjKv7Wnlwi6D+sawbZA/i8aEwzpgoLi54BW2ql8bF
ZVSsnk2cqOwNRs77nuJTlgY+W8dbNWhYio4Tj8O5zr9eu0w66OCjCCvdtuTYozfB+WVK1U/gC9Hk
VIBHGcDRIcku1vC/s/G7/IrJ7SrMRAgHYZMUXcviqKEFAgitCpceWKv/x9TiWnh2/flFIAjjaOZM
1IkCCDWxWgCNdMplioaEdU/LjOVAqEItzA+tFMV/uiBwQZQ3ly7PXAi7ISjx+FT1HQ55mjSt05F5
/e+ykkewloePrQ/ZcqTCgU2lUJOifZCyXpVUfcvaS05AAncy72+kd6GofrecyoAVkvhB5HbJKnzE
KGP/IL+xWJSwFpeAeWUrllWtPHkgGpBVsGqUNZ3ixzREsgu/wS1+0fRHqY6DJVgF/9VXuX4YF/gy
2giy791mYl0G4R2jLiSCrdqJOnxMtD3eVfeMHAiS6IW0+jQI4XRPpUIE9NHea+tOv5h9KNmWxEv1
FL+sUcgrdhYi53INrAwch5FuTpMRALShxUCHXkA+g88VeQ2sIGJffHLGZuXb7nwKsEU7jqGR5GC2
j9d7WQB6TET/vpPozDMxRB0b9ucq3RrewRQAVVR0IHI1OCXTguNjUXB0Kr29PqrGKpFutwipfmct
D7gqiWIVo3tXmBYn1Itg0yQFsJMn/wDtvpW3ONwUuM4BcDACC1wWeEaJr1BqKEamUla0WF3YD3QX
3dKIyV+ue0PIfKFxshgoXL7FYtcyQJqX1f+f8WbG/KHgtTxnokyySm849zbxwQk6jDp7rB/u9kCa
btEEtHirbWoDuGLAy0syA7f/7LVZ+17IC2OZ3W1EMlinCgyOL7b1ih+SZSH4XxWYRTuJb41nJe/K
nqDd46IZS6hAOrP8hYinlVPzEGkF6BAJRyz9/TG9ML90+fKr+PjlYKm3oedxkKAsv4GhWHxsQyuF
0iGNOgpOmIjeZHyZM8+ax130hCoDv0mJILC3cFOx4l7uw1uwa/2Hgc9diQrSkVEJExjhtKpJSd5Y
nYHAaf3zwykRr5xpkA1eF5UFDbDiHth6UNyC4gYN0Y0biTDXS4gIau6Z91kwUJoch8v0o4Bt2ANa
wdTj+Zpk078GNklezi5mwKLV4w+f2Ba1ZQs9JePhc43JdG/8JPs08IWm9XxBOAQVNnrC4UKBS2AQ
cJc59JjB2VDyEH67J0jqTya5d05nDqbos3r4KjVpXu1FxhBZv2iBLexm+ZgRb/ZeY+C6k7S1sl0W
dkpPbHNYtkZLbRy/hPHa1IbqsAK7G3AI6xBmyWNf/1IYN84DHrXlaW75UQtaHnWVaoHLI1wEGqXB
k+P+1LjAI9HNvdOXZn98wzqtW1o+K8pnULE9g2NzD4jslt30zM4r/RitK1S0njuEOgI58ST2DEXq
LUaL/epAxRmLWDmSSWpnofZ0kltFmbOLy+gtS3q8Cdx1vcROO5la24lybM2G9/14Tki3CuNx5J0Z
nEctilV1zhcCMKylgbOyeFQoqH+pZCUYK78R/CkARSr2ikSYtQ4ZtSdNnP94D/ce7wXLHDPpRcbI
xPudXgFLRHShMNikwgD6dRJm6juuY3oUxI0DtN9feiNnbvQtwHpchKTGo721kq27Bt9pRDWFsMi4
8O0DntBJial+VX4Vu4bNf0LmkcEGeyFS7LjILZJr1kvVMX95BBpYgQEmTWWAf/lBItTo76mCXSdk
OLUK81lS9lXco5QoS0nSyRfdFhBgcNbQaAIxPTzxZuRLZIjpODkZOftmp93GWbKZJjIqXhOarSAX
XeRr7efz+56u7SX00bh5utOnRDylPywcZdTthXJToOkLfn7YvOOti2lystrvASjY/FyAb+6ciRug
HEJZHRY17rCBKUTWtX7nvgx7SWnAFTJjqldFlGwvRO90Nztjt6cGOjOG5GVP+FBNfErAXaxsGHLl
cfjPqU+NC93Kdj+PFeYgfA0VQcZd5ci7c1Dj6R/n2QPnYfk7kVr+nu1xecJ/VFD3IrLWS886M3Hx
BoBd6rGz+FuO+h/ydSRxSwhTcjPnTnDSFk4//1tmh0x3pNj09FN0AoV8FMbVl8jos577+8jI2kw0
cszz84RSiNSfs17qjqKWhNNg+txnMINqlB3pphVlYvpR5vAX/IGFWx5KWoU13Pw2ZyFQYRNngmAj
LyjJ7XrY8tcnF2O+w9VbzKbDWxwnFwNTrnv/wT+L+Y7ozgwocFPSbJFZwYZBsjbMrdo57Bdax1/j
T1XHyIMDoYbxPgCn0b6Mnwy2roDLhe6uKF2/NEIG7cxM4zjuW8pI7YpoZSZwlKGb9HEGyWRmzmmR
030ne0atwA5xnBc7sK38LHRFDk7btG7kSnwyQm+zuI8a1NPDRdNXwJ6t3AXsAARhvB0iUkFkkVOG
GpKF3a9C2ug+SsghOJ6d1LJ8hOrALQIuTSyzB84vsvi0pzNs1MYJfAIQa4C+n8wlB+0TCrdOylxi
ZMam0/wr3MIx/3Qaot8MZLRMfmnTrSuQy28eJseZb9QdOccwaw5a4NZLmjig4+vgWJ+6GsQk3hj/
LPBSg0N7SlNgWekxfbHO05Mc+GmSN3tcYv4+9jckhvuYdAsFIvCFQgO46DQ9oWNPQWkiDqlDY9OP
NCZiZWOrzMVPN8zV2KmBmqBNSSvWasHxld0K4xQR8EenPDSSGHP9wo07nA77i7l92EDGaBTi1f9y
sH/2FkXOSpDTVrljR48fAwouG+BS3hPMK//qDrrMXxB4tfvSl+BQoCuAdepXTAfXduyKrFB5zYsr
+n1Uv/JPMWwnl5VLczQ3aHkh19JcQhiCjGS6vxcJHzfc+aILyr7gKb2ubSouIsY0yc8g6IYOnoDD
+XCRuEPOag4IRbv1WsC1IXyDe1Twpr/0LemGmUMcjsHh5HV21zwl5x/lcOGi32Fr+x8uaXsEGicO
XSUvCuZCHSwT6P+cUiF0+l9yHyUMuZkJ5bji5Yld9aeQxNZpstPbDvl2A5SKfc1ohsLoIhq4i3ds
40Y8d7i2Lp4CiaG9hkXTPB1AAliZYPbUTICsrZYRQRTfGmJPIVFJvjrwJI6d5RDugowkaju8AoYM
A+qMd8H7lDfq/rtnVrPKfufESxkB1Q2ALqFXbmTwcM+58yiiuwOnm5+smLvQeFigyRO2VLRMt3/v
okt0PssCTyHWuQVNRTYGBWIoWTP9yM/WoQ2TN8mtfQ6JGUQcLUBIWY1pBc69WwCe4DkHCYeMRemX
I3yjba++DukMOBoNHicuBVSJ3zGu/z9/H7OhZ+oGkD13SpqqaUHIs2tqA6Oyvueq93lu3TpZJdDv
GeW0anTk6kyZhgAR/SFN/B+FMXyCZQsCVkzaZCYphsEwLeJcCOJWbeXlQJHkGhz1v6wzyyJpYxOJ
5ZByyfsgjFVaX+ti9t3wtSTYvgwOtAvLkhY4/lH7AtUYOgQS4VODERXgQyDNdlao1BxfucBDptKr
JOBgh5wzCh5YE74cGHFt6qhO2G5PK/sFnu1/ChKyItuC4UMANJ6QAqYIYJG41vEatfbhLqSUQykk
W6UWgOe7wq/mR6g8FdKbsi794gzePbNtqgirBr7d98iPjyP3wzJyKwSeuK+Ul+9SCPGZDt2iOAqe
1abCmPHPKZAWV0fVlom0I8suA5RE4X9n8cONRIvwdXUW2rz8ritgIXw8dKY6fH7YW+OuU+zdJ1Pn
k5ZkILe76niAZTy7g5njgCP1EheRDDBOF9k/SSMgolMK/Po3l/JNMxtqmtuGLEOQvAaTpl5U9Wpc
cXaBUTC0+Bqscug/H8slnlhAFiraXuhaP2Ie+ePRklYXTXFJvK3AfsLgKWBMXVz2xQd4BW0uIIBV
TWj+JF2fqemnzLEg0d5NL6L5QbFTbGkJ74866G7oPoCn0JLELYBsfzKEGoRfsizpey6DACxHhiau
GoKpAFHGTrZIrJV/Kx515VpHs9sgP2C7qekxyz1qBJOAv4ZLtoKATp1I/IWYBueneWy2NcLJnyOE
GmrQvtBcvQ+Zt6iyeaBCmCV0a2CLtXSSgxvJwKgNU451EokkyXZRIhcY7a7Td6IFE032YZiezEiL
pXKv2TjIxIfmwp9EmgXwVKbddXaIzwYrL2B8bmw3sbAc2xHBLN6h2tc6Os53UshsA2CdkgV47ah1
NbUNm/VAZr0cH14X9pxpOWwqfzO9tf/cl88huNRqhgcteFoLHUPUlQmZQusdl3gO7s/d6etSencj
EoUBlUluaUAQtOEzHNCn7ea2UbOlSItHMDTVo/+LQpqWwLwQU75oN5AhQunjfB/WcQf8n3Mrg0oY
baOKUPd5QXTMkjfZsoRQ59VuyTGhMwB4MDva2c0vIWGplhxDdB2IkHVyqzr3fX9Jw/eO08X/Ir2E
U5eukT/g+ho//dCCk/Q6WlCYqVh5Lm8/rHcIXmEKt1gE+VMO7GmzZ2Eb6hmkHq5neZKfpHJPCU2v
rbBEzJYG84dAASLk/UgQIkKjGcmT9LoE0irT0NtRK6Qr1YGOnasI
`protect end_protected
